module dft_testbench();

initial begin 
	$dumpfile("fft_fx64_it_rdx8_w512.vcd");
	$dumpvars(4);
end

   reg clk, reset, next;
   wire next_out;
   integer i, j, k, l, m;
   reg [15:0] counter;
   reg [63:0] in [1023:0];
   wire [63:0] X0;
   wire [63:0] Y0;
   wire [63:0] X1;
   wire [63:0] Y1;
   wire [63:0] X2;
   wire [63:0] Y2;
   wire [63:0] X3;
   wire [63:0] Y3;
   wire [63:0] X4;
   wire [63:0] Y4;
   wire [63:0] X5;
   wire [63:0] Y5;
   wire [63:0] X6;
   wire [63:0] Y6;
   wire [63:0] X7;
   wire [63:0] Y7;
   wire [63:0] X8;
   wire [63:0] Y8;
   wire [63:0] X9;
   wire [63:0] Y9;
   wire [63:0] X10;
   wire [63:0] Y10;
   wire [63:0] X11;
   wire [63:0] Y11;
   wire [63:0] X12;
   wire [63:0] Y12;
   wire [63:0] X13;
   wire [63:0] Y13;
   wire [63:0] X14;
   wire [63:0] Y14;
   wire [63:0] X15;
   wire [63:0] Y15;
   wire [63:0] X16;
   wire [63:0] Y16;
   wire [63:0] X17;
   wire [63:0] Y17;
   wire [63:0] X18;
   wire [63:0] Y18;
   wire [63:0] X19;
   wire [63:0] Y19;
   wire [63:0] X20;
   wire [63:0] Y20;
   wire [63:0] X21;
   wire [63:0] Y21;
   wire [63:0] X22;
   wire [63:0] Y22;
   wire [63:0] X23;
   wire [63:0] Y23;
   wire [63:0] X24;
   wire [63:0] Y24;
   wire [63:0] X25;
   wire [63:0] Y25;
   wire [63:0] X26;
   wire [63:0] Y26;
   wire [63:0] X27;
   wire [63:0] Y27;
   wire [63:0] X28;
   wire [63:0] Y28;
   wire [63:0] X29;
   wire [63:0] Y29;
   wire [63:0] X30;
   wire [63:0] Y30;
   wire [63:0] X31;
   wire [63:0] Y31;
   wire [63:0] X32;
   wire [63:0] Y32;
   wire [63:0] X33;
   wire [63:0] Y33;
   wire [63:0] X34;
   wire [63:0] Y34;
   wire [63:0] X35;
   wire [63:0] Y35;
   wire [63:0] X36;
   wire [63:0] Y36;
   wire [63:0] X37;
   wire [63:0] Y37;
   wire [63:0] X38;
   wire [63:0] Y38;
   wire [63:0] X39;
   wire [63:0] Y39;
   wire [63:0] X40;
   wire [63:0] Y40;
   wire [63:0] X41;
   wire [63:0] Y41;
   wire [63:0] X42;
   wire [63:0] Y42;
   wire [63:0] X43;
   wire [63:0] Y43;
   wire [63:0] X44;
   wire [63:0] Y44;
   wire [63:0] X45;
   wire [63:0] Y45;
   wire [63:0] X46;
   wire [63:0] Y46;
   wire [63:0] X47;
   wire [63:0] Y47;
   wire [63:0] X48;
   wire [63:0] Y48;
   wire [63:0] X49;
   wire [63:0] Y49;
   wire [63:0] X50;
   wire [63:0] Y50;
   wire [63:0] X51;
   wire [63:0] Y51;
   wire [63:0] X52;
   wire [63:0] Y52;
   wire [63:0] X53;
   wire [63:0] Y53;
   wire [63:0] X54;
   wire [63:0] Y54;
   wire [63:0] X55;
   wire [63:0] Y55;
   wire [63:0] X56;
   wire [63:0] Y56;
   wire [63:0] X57;
   wire [63:0] Y57;
   wire [63:0] X58;
   wire [63:0] Y58;
   wire [63:0] X59;
   wire [63:0] Y59;
   wire [63:0] X60;
   wire [63:0] Y60;
   wire [63:0] X61;
   wire [63:0] Y61;
   wire [63:0] X62;
   wire [63:0] Y62;
   wire [63:0] X63;
   wire [63:0] Y63;
   wire [63:0] X64;
   wire [63:0] Y64;
   wire [63:0] X65;
   wire [63:0] Y65;
   wire [63:0] X66;
   wire [63:0] Y66;
   wire [63:0] X67;
   wire [63:0] Y67;
   wire [63:0] X68;
   wire [63:0] Y68;
   wire [63:0] X69;
   wire [63:0] Y69;
   wire [63:0] X70;
   wire [63:0] Y70;
   wire [63:0] X71;
   wire [63:0] Y71;
   wire [63:0] X72;
   wire [63:0] Y72;
   wire [63:0] X73;
   wire [63:0] Y73;
   wire [63:0] X74;
   wire [63:0] Y74;
   wire [63:0] X75;
   wire [63:0] Y75;
   wire [63:0] X76;
   wire [63:0] Y76;
   wire [63:0] X77;
   wire [63:0] Y77;
   wire [63:0] X78;
   wire [63:0] Y78;
   wire [63:0] X79;
   wire [63:0] Y79;
   wire [63:0] X80;
   wire [63:0] Y80;
   wire [63:0] X81;
   wire [63:0] Y81;
   wire [63:0] X82;
   wire [63:0] Y82;
   wire [63:0] X83;
   wire [63:0] Y83;
   wire [63:0] X84;
   wire [63:0] Y84;
   wire [63:0] X85;
   wire [63:0] Y85;
   wire [63:0] X86;
   wire [63:0] Y86;
   wire [63:0] X87;
   wire [63:0] Y87;
   wire [63:0] X88;
   wire [63:0] Y88;
   wire [63:0] X89;
   wire [63:0] Y89;
   wire [63:0] X90;
   wire [63:0] Y90;
   wire [63:0] X91;
   wire [63:0] Y91;
   wire [63:0] X92;
   wire [63:0] Y92;
   wire [63:0] X93;
   wire [63:0] Y93;
   wire [63:0] X94;
   wire [63:0] Y94;
   wire [63:0] X95;
   wire [63:0] Y95;
   wire [63:0] X96;
   wire [63:0] Y96;
   wire [63:0] X97;
   wire [63:0] Y97;
   wire [63:0] X98;
   wire [63:0] Y98;
   wire [63:0] X99;
   wire [63:0] Y99;
   wire [63:0] X100;
   wire [63:0] Y100;
   wire [63:0] X101;
   wire [63:0] Y101;
   wire [63:0] X102;
   wire [63:0] Y102;
   wire [63:0] X103;
   wire [63:0] Y103;
   wire [63:0] X104;
   wire [63:0] Y104;
   wire [63:0] X105;
   wire [63:0] Y105;
   wire [63:0] X106;
   wire [63:0] Y106;
   wire [63:0] X107;
   wire [63:0] Y107;
   wire [63:0] X108;
   wire [63:0] Y108;
   wire [63:0] X109;
   wire [63:0] Y109;
   wire [63:0] X110;
   wire [63:0] Y110;
   wire [63:0] X111;
   wire [63:0] Y111;
   wire [63:0] X112;
   wire [63:0] Y112;
   wire [63:0] X113;
   wire [63:0] Y113;
   wire [63:0] X114;
   wire [63:0] Y114;
   wire [63:0] X115;
   wire [63:0] Y115;
   wire [63:0] X116;
   wire [63:0] Y116;
   wire [63:0] X117;
   wire [63:0] Y117;
   wire [63:0] X118;
   wire [63:0] Y118;
   wire [63:0] X119;
   wire [63:0] Y119;
   wire [63:0] X120;
   wire [63:0] Y120;
   wire [63:0] X121;
   wire [63:0] Y121;
   wire [63:0] X122;
   wire [63:0] Y122;
   wire [63:0] X123;
   wire [63:0] Y123;
   wire [63:0] X124;
   wire [63:0] Y124;
   wire [63:0] X125;
   wire [63:0] Y125;
   wire [63:0] X126;
   wire [63:0] Y126;
   wire [63:0] X127;
   wire [63:0] Y127;
   wire [63:0] X128;
   wire [63:0] Y128;
   wire [63:0] X129;
   wire [63:0] Y129;
   wire [63:0] X130;
   wire [63:0] Y130;
   wire [63:0] X131;
   wire [63:0] Y131;
   wire [63:0] X132;
   wire [63:0] Y132;
   wire [63:0] X133;
   wire [63:0] Y133;
   wire [63:0] X134;
   wire [63:0] Y134;
   wire [63:0] X135;
   wire [63:0] Y135;
   wire [63:0] X136;
   wire [63:0] Y136;
   wire [63:0] X137;
   wire [63:0] Y137;
   wire [63:0] X138;
   wire [63:0] Y138;
   wire [63:0] X139;
   wire [63:0] Y139;
   wire [63:0] X140;
   wire [63:0] Y140;
   wire [63:0] X141;
   wire [63:0] Y141;
   wire [63:0] X142;
   wire [63:0] Y142;
   wire [63:0] X143;
   wire [63:0] Y143;
   wire [63:0] X144;
   wire [63:0] Y144;
   wire [63:0] X145;
   wire [63:0] Y145;
   wire [63:0] X146;
   wire [63:0] Y146;
   wire [63:0] X147;
   wire [63:0] Y147;
   wire [63:0] X148;
   wire [63:0] Y148;
   wire [63:0] X149;
   wire [63:0] Y149;
   wire [63:0] X150;
   wire [63:0] Y150;
   wire [63:0] X151;
   wire [63:0] Y151;
   wire [63:0] X152;
   wire [63:0] Y152;
   wire [63:0] X153;
   wire [63:0] Y153;
   wire [63:0] X154;
   wire [63:0] Y154;
   wire [63:0] X155;
   wire [63:0] Y155;
   wire [63:0] X156;
   wire [63:0] Y156;
   wire [63:0] X157;
   wire [63:0] Y157;
   wire [63:0] X158;
   wire [63:0] Y158;
   wire [63:0] X159;
   wire [63:0] Y159;
   wire [63:0] X160;
   wire [63:0] Y160;
   wire [63:0] X161;
   wire [63:0] Y161;
   wire [63:0] X162;
   wire [63:0] Y162;
   wire [63:0] X163;
   wire [63:0] Y163;
   wire [63:0] X164;
   wire [63:0] Y164;
   wire [63:0] X165;
   wire [63:0] Y165;
   wire [63:0] X166;
   wire [63:0] Y166;
   wire [63:0] X167;
   wire [63:0] Y167;
   wire [63:0] X168;
   wire [63:0] Y168;
   wire [63:0] X169;
   wire [63:0] Y169;
   wire [63:0] X170;
   wire [63:0] Y170;
   wire [63:0] X171;
   wire [63:0] Y171;
   wire [63:0] X172;
   wire [63:0] Y172;
   wire [63:0] X173;
   wire [63:0] Y173;
   wire [63:0] X174;
   wire [63:0] Y174;
   wire [63:0] X175;
   wire [63:0] Y175;
   wire [63:0] X176;
   wire [63:0] Y176;
   wire [63:0] X177;
   wire [63:0] Y177;
   wire [63:0] X178;
   wire [63:0] Y178;
   wire [63:0] X179;
   wire [63:0] Y179;
   wire [63:0] X180;
   wire [63:0] Y180;
   wire [63:0] X181;
   wire [63:0] Y181;
   wire [63:0] X182;
   wire [63:0] Y182;
   wire [63:0] X183;
   wire [63:0] Y183;
   wire [63:0] X184;
   wire [63:0] Y184;
   wire [63:0] X185;
   wire [63:0] Y185;
   wire [63:0] X186;
   wire [63:0] Y186;
   wire [63:0] X187;
   wire [63:0] Y187;
   wire [63:0] X188;
   wire [63:0] Y188;
   wire [63:0] X189;
   wire [63:0] Y189;
   wire [63:0] X190;
   wire [63:0] Y190;
   wire [63:0] X191;
   wire [63:0] Y191;
   wire [63:0] X192;
   wire [63:0] Y192;
   wire [63:0] X193;
   wire [63:0] Y193;
   wire [63:0] X194;
   wire [63:0] Y194;
   wire [63:0] X195;
   wire [63:0] Y195;
   wire [63:0] X196;
   wire [63:0] Y196;
   wire [63:0] X197;
   wire [63:0] Y197;
   wire [63:0] X198;
   wire [63:0] Y198;
   wire [63:0] X199;
   wire [63:0] Y199;
   wire [63:0] X200;
   wire [63:0] Y200;
   wire [63:0] X201;
   wire [63:0] Y201;
   wire [63:0] X202;
   wire [63:0] Y202;
   wire [63:0] X203;
   wire [63:0] Y203;
   wire [63:0] X204;
   wire [63:0] Y204;
   wire [63:0] X205;
   wire [63:0] Y205;
   wire [63:0] X206;
   wire [63:0] Y206;
   wire [63:0] X207;
   wire [63:0] Y207;
   wire [63:0] X208;
   wire [63:0] Y208;
   wire [63:0] X209;
   wire [63:0] Y209;
   wire [63:0] X210;
   wire [63:0] Y210;
   wire [63:0] X211;
   wire [63:0] Y211;
   wire [63:0] X212;
   wire [63:0] Y212;
   wire [63:0] X213;
   wire [63:0] Y213;
   wire [63:0] X214;
   wire [63:0] Y214;
   wire [63:0] X215;
   wire [63:0] Y215;
   wire [63:0] X216;
   wire [63:0] Y216;
   wire [63:0] X217;
   wire [63:0] Y217;
   wire [63:0] X218;
   wire [63:0] Y218;
   wire [63:0] X219;
   wire [63:0] Y219;
   wire [63:0] X220;
   wire [63:0] Y220;
   wire [63:0] X221;
   wire [63:0] Y221;
   wire [63:0] X222;
   wire [63:0] Y222;
   wire [63:0] X223;
   wire [63:0] Y223;
   wire [63:0] X224;
   wire [63:0] Y224;
   wire [63:0] X225;
   wire [63:0] Y225;
   wire [63:0] X226;
   wire [63:0] Y226;
   wire [63:0] X227;
   wire [63:0] Y227;
   wire [63:0] X228;
   wire [63:0] Y228;
   wire [63:0] X229;
   wire [63:0] Y229;
   wire [63:0] X230;
   wire [63:0] Y230;
   wire [63:0] X231;
   wire [63:0] Y231;
   wire [63:0] X232;
   wire [63:0] Y232;
   wire [63:0] X233;
   wire [63:0] Y233;
   wire [63:0] X234;
   wire [63:0] Y234;
   wire [63:0] X235;
   wire [63:0] Y235;
   wire [63:0] X236;
   wire [63:0] Y236;
   wire [63:0] X237;
   wire [63:0] Y237;
   wire [63:0] X238;
   wire [63:0] Y238;
   wire [63:0] X239;
   wire [63:0] Y239;
   wire [63:0] X240;
   wire [63:0] Y240;
   wire [63:0] X241;
   wire [63:0] Y241;
   wire [63:0] X242;
   wire [63:0] Y242;
   wire [63:0] X243;
   wire [63:0] Y243;
   wire [63:0] X244;
   wire [63:0] Y244;
   wire [63:0] X245;
   wire [63:0] Y245;
   wire [63:0] X246;
   wire [63:0] Y246;
   wire [63:0] X247;
   wire [63:0] Y247;
   wire [63:0] X248;
   wire [63:0] Y248;
   wire [63:0] X249;
   wire [63:0] Y249;
   wire [63:0] X250;
   wire [63:0] Y250;
   wire [63:0] X251;
   wire [63:0] Y251;
   wire [63:0] X252;
   wire [63:0] Y252;
   wire [63:0] X253;
   wire [63:0] Y253;
   wire [63:0] X254;
   wire [63:0] Y254;
   wire [63:0] X255;
   wire [63:0] Y255;
   wire [63:0] X256;
   wire [63:0] Y256;
   wire [63:0] X257;
   wire [63:0] Y257;
   wire [63:0] X258;
   wire [63:0] Y258;
   wire [63:0] X259;
   wire [63:0] Y259;
   wire [63:0] X260;
   wire [63:0] Y260;
   wire [63:0] X261;
   wire [63:0] Y261;
   wire [63:0] X262;
   wire [63:0] Y262;
   wire [63:0] X263;
   wire [63:0] Y263;
   wire [63:0] X264;
   wire [63:0] Y264;
   wire [63:0] X265;
   wire [63:0] Y265;
   wire [63:0] X266;
   wire [63:0] Y266;
   wire [63:0] X267;
   wire [63:0] Y267;
   wire [63:0] X268;
   wire [63:0] Y268;
   wire [63:0] X269;
   wire [63:0] Y269;
   wire [63:0] X270;
   wire [63:0] Y270;
   wire [63:0] X271;
   wire [63:0] Y271;
   wire [63:0] X272;
   wire [63:0] Y272;
   wire [63:0] X273;
   wire [63:0] Y273;
   wire [63:0] X274;
   wire [63:0] Y274;
   wire [63:0] X275;
   wire [63:0] Y275;
   wire [63:0] X276;
   wire [63:0] Y276;
   wire [63:0] X277;
   wire [63:0] Y277;
   wire [63:0] X278;
   wire [63:0] Y278;
   wire [63:0] X279;
   wire [63:0] Y279;
   wire [63:0] X280;
   wire [63:0] Y280;
   wire [63:0] X281;
   wire [63:0] Y281;
   wire [63:0] X282;
   wire [63:0] Y282;
   wire [63:0] X283;
   wire [63:0] Y283;
   wire [63:0] X284;
   wire [63:0] Y284;
   wire [63:0] X285;
   wire [63:0] Y285;
   wire [63:0] X286;
   wire [63:0] Y286;
   wire [63:0] X287;
   wire [63:0] Y287;
   wire [63:0] X288;
   wire [63:0] Y288;
   wire [63:0] X289;
   wire [63:0] Y289;
   wire [63:0] X290;
   wire [63:0] Y290;
   wire [63:0] X291;
   wire [63:0] Y291;
   wire [63:0] X292;
   wire [63:0] Y292;
   wire [63:0] X293;
   wire [63:0] Y293;
   wire [63:0] X294;
   wire [63:0] Y294;
   wire [63:0] X295;
   wire [63:0] Y295;
   wire [63:0] X296;
   wire [63:0] Y296;
   wire [63:0] X297;
   wire [63:0] Y297;
   wire [63:0] X298;
   wire [63:0] Y298;
   wire [63:0] X299;
   wire [63:0] Y299;
   wire [63:0] X300;
   wire [63:0] Y300;
   wire [63:0] X301;
   wire [63:0] Y301;
   wire [63:0] X302;
   wire [63:0] Y302;
   wire [63:0] X303;
   wire [63:0] Y303;
   wire [63:0] X304;
   wire [63:0] Y304;
   wire [63:0] X305;
   wire [63:0] Y305;
   wire [63:0] X306;
   wire [63:0] Y306;
   wire [63:0] X307;
   wire [63:0] Y307;
   wire [63:0] X308;
   wire [63:0] Y308;
   wire [63:0] X309;
   wire [63:0] Y309;
   wire [63:0] X310;
   wire [63:0] Y310;
   wire [63:0] X311;
   wire [63:0] Y311;
   wire [63:0] X312;
   wire [63:0] Y312;
   wire [63:0] X313;
   wire [63:0] Y313;
   wire [63:0] X314;
   wire [63:0] Y314;
   wire [63:0] X315;
   wire [63:0] Y315;
   wire [63:0] X316;
   wire [63:0] Y316;
   wire [63:0] X317;
   wire [63:0] Y317;
   wire [63:0] X318;
   wire [63:0] Y318;
   wire [63:0] X319;
   wire [63:0] Y319;
   wire [63:0] X320;
   wire [63:0] Y320;
   wire [63:0] X321;
   wire [63:0] Y321;
   wire [63:0] X322;
   wire [63:0] Y322;
   wire [63:0] X323;
   wire [63:0] Y323;
   wire [63:0] X324;
   wire [63:0] Y324;
   wire [63:0] X325;
   wire [63:0] Y325;
   wire [63:0] X326;
   wire [63:0] Y326;
   wire [63:0] X327;
   wire [63:0] Y327;
   wire [63:0] X328;
   wire [63:0] Y328;
   wire [63:0] X329;
   wire [63:0] Y329;
   wire [63:0] X330;
   wire [63:0] Y330;
   wire [63:0] X331;
   wire [63:0] Y331;
   wire [63:0] X332;
   wire [63:0] Y332;
   wire [63:0] X333;
   wire [63:0] Y333;
   wire [63:0] X334;
   wire [63:0] Y334;
   wire [63:0] X335;
   wire [63:0] Y335;
   wire [63:0] X336;
   wire [63:0] Y336;
   wire [63:0] X337;
   wire [63:0] Y337;
   wire [63:0] X338;
   wire [63:0] Y338;
   wire [63:0] X339;
   wire [63:0] Y339;
   wire [63:0] X340;
   wire [63:0] Y340;
   wire [63:0] X341;
   wire [63:0] Y341;
   wire [63:0] X342;
   wire [63:0] Y342;
   wire [63:0] X343;
   wire [63:0] Y343;
   wire [63:0] X344;
   wire [63:0] Y344;
   wire [63:0] X345;
   wire [63:0] Y345;
   wire [63:0] X346;
   wire [63:0] Y346;
   wire [63:0] X347;
   wire [63:0] Y347;
   wire [63:0] X348;
   wire [63:0] Y348;
   wire [63:0] X349;
   wire [63:0] Y349;
   wire [63:0] X350;
   wire [63:0] Y350;
   wire [63:0] X351;
   wire [63:0] Y351;
   wire [63:0] X352;
   wire [63:0] Y352;
   wire [63:0] X353;
   wire [63:0] Y353;
   wire [63:0] X354;
   wire [63:0] Y354;
   wire [63:0] X355;
   wire [63:0] Y355;
   wire [63:0] X356;
   wire [63:0] Y356;
   wire [63:0] X357;
   wire [63:0] Y357;
   wire [63:0] X358;
   wire [63:0] Y358;
   wire [63:0] X359;
   wire [63:0] Y359;
   wire [63:0] X360;
   wire [63:0] Y360;
   wire [63:0] X361;
   wire [63:0] Y361;
   wire [63:0] X362;
   wire [63:0] Y362;
   wire [63:0] X363;
   wire [63:0] Y363;
   wire [63:0] X364;
   wire [63:0] Y364;
   wire [63:0] X365;
   wire [63:0] Y365;
   wire [63:0] X366;
   wire [63:0] Y366;
   wire [63:0] X367;
   wire [63:0] Y367;
   wire [63:0] X368;
   wire [63:0] Y368;
   wire [63:0] X369;
   wire [63:0] Y369;
   wire [63:0] X370;
   wire [63:0] Y370;
   wire [63:0] X371;
   wire [63:0] Y371;
   wire [63:0] X372;
   wire [63:0] Y372;
   wire [63:0] X373;
   wire [63:0] Y373;
   wire [63:0] X374;
   wire [63:0] Y374;
   wire [63:0] X375;
   wire [63:0] Y375;
   wire [63:0] X376;
   wire [63:0] Y376;
   wire [63:0] X377;
   wire [63:0] Y377;
   wire [63:0] X378;
   wire [63:0] Y378;
   wire [63:0] X379;
   wire [63:0] Y379;
   wire [63:0] X380;
   wire [63:0] Y380;
   wire [63:0] X381;
   wire [63:0] Y381;
   wire [63:0] X382;
   wire [63:0] Y382;
   wire [63:0] X383;
   wire [63:0] Y383;
   wire [63:0] X384;
   wire [63:0] Y384;
   wire [63:0] X385;
   wire [63:0] Y385;
   wire [63:0] X386;
   wire [63:0] Y386;
   wire [63:0] X387;
   wire [63:0] Y387;
   wire [63:0] X388;
   wire [63:0] Y388;
   wire [63:0] X389;
   wire [63:0] Y389;
   wire [63:0] X390;
   wire [63:0] Y390;
   wire [63:0] X391;
   wire [63:0] Y391;
   wire [63:0] X392;
   wire [63:0] Y392;
   wire [63:0] X393;
   wire [63:0] Y393;
   wire [63:0] X394;
   wire [63:0] Y394;
   wire [63:0] X395;
   wire [63:0] Y395;
   wire [63:0] X396;
   wire [63:0] Y396;
   wire [63:0] X397;
   wire [63:0] Y397;
   wire [63:0] X398;
   wire [63:0] Y398;
   wire [63:0] X399;
   wire [63:0] Y399;
   wire [63:0] X400;
   wire [63:0] Y400;
   wire [63:0] X401;
   wire [63:0] Y401;
   wire [63:0] X402;
   wire [63:0] Y402;
   wire [63:0] X403;
   wire [63:0] Y403;
   wire [63:0] X404;
   wire [63:0] Y404;
   wire [63:0] X405;
   wire [63:0] Y405;
   wire [63:0] X406;
   wire [63:0] Y406;
   wire [63:0] X407;
   wire [63:0] Y407;
   wire [63:0] X408;
   wire [63:0] Y408;
   wire [63:0] X409;
   wire [63:0] Y409;
   wire [63:0] X410;
   wire [63:0] Y410;
   wire [63:0] X411;
   wire [63:0] Y411;
   wire [63:0] X412;
   wire [63:0] Y412;
   wire [63:0] X413;
   wire [63:0] Y413;
   wire [63:0] X414;
   wire [63:0] Y414;
   wire [63:0] X415;
   wire [63:0] Y415;
   wire [63:0] X416;
   wire [63:0] Y416;
   wire [63:0] X417;
   wire [63:0] Y417;
   wire [63:0] X418;
   wire [63:0] Y418;
   wire [63:0] X419;
   wire [63:0] Y419;
   wire [63:0] X420;
   wire [63:0] Y420;
   wire [63:0] X421;
   wire [63:0] Y421;
   wire [63:0] X422;
   wire [63:0] Y422;
   wire [63:0] X423;
   wire [63:0] Y423;
   wire [63:0] X424;
   wire [63:0] Y424;
   wire [63:0] X425;
   wire [63:0] Y425;
   wire [63:0] X426;
   wire [63:0] Y426;
   wire [63:0] X427;
   wire [63:0] Y427;
   wire [63:0] X428;
   wire [63:0] Y428;
   wire [63:0] X429;
   wire [63:0] Y429;
   wire [63:0] X430;
   wire [63:0] Y430;
   wire [63:0] X431;
   wire [63:0] Y431;
   wire [63:0] X432;
   wire [63:0] Y432;
   wire [63:0] X433;
   wire [63:0] Y433;
   wire [63:0] X434;
   wire [63:0] Y434;
   wire [63:0] X435;
   wire [63:0] Y435;
   wire [63:0] X436;
   wire [63:0] Y436;
   wire [63:0] X437;
   wire [63:0] Y437;
   wire [63:0] X438;
   wire [63:0] Y438;
   wire [63:0] X439;
   wire [63:0] Y439;
   wire [63:0] X440;
   wire [63:0] Y440;
   wire [63:0] X441;
   wire [63:0] Y441;
   wire [63:0] X442;
   wire [63:0] Y442;
   wire [63:0] X443;
   wire [63:0] Y443;
   wire [63:0] X444;
   wire [63:0] Y444;
   wire [63:0] X445;
   wire [63:0] Y445;
   wire [63:0] X446;
   wire [63:0] Y446;
   wire [63:0] X447;
   wire [63:0] Y447;
   wire [63:0] X448;
   wire [63:0] Y448;
   wire [63:0] X449;
   wire [63:0] Y449;
   wire [63:0] X450;
   wire [63:0] Y450;
   wire [63:0] X451;
   wire [63:0] Y451;
   wire [63:0] X452;
   wire [63:0] Y452;
   wire [63:0] X453;
   wire [63:0] Y453;
   wire [63:0] X454;
   wire [63:0] Y454;
   wire [63:0] X455;
   wire [63:0] Y455;
   wire [63:0] X456;
   wire [63:0] Y456;
   wire [63:0] X457;
   wire [63:0] Y457;
   wire [63:0] X458;
   wire [63:0] Y458;
   wire [63:0] X459;
   wire [63:0] Y459;
   wire [63:0] X460;
   wire [63:0] Y460;
   wire [63:0] X461;
   wire [63:0] Y461;
   wire [63:0] X462;
   wire [63:0] Y462;
   wire [63:0] X463;
   wire [63:0] Y463;
   wire [63:0] X464;
   wire [63:0] Y464;
   wire [63:0] X465;
   wire [63:0] Y465;
   wire [63:0] X466;
   wire [63:0] Y466;
   wire [63:0] X467;
   wire [63:0] Y467;
   wire [63:0] X468;
   wire [63:0] Y468;
   wire [63:0] X469;
   wire [63:0] Y469;
   wire [63:0] X470;
   wire [63:0] Y470;
   wire [63:0] X471;
   wire [63:0] Y471;
   wire [63:0] X472;
   wire [63:0] Y472;
   wire [63:0] X473;
   wire [63:0] Y473;
   wire [63:0] X474;
   wire [63:0] Y474;
   wire [63:0] X475;
   wire [63:0] Y475;
   wire [63:0] X476;
   wire [63:0] Y476;
   wire [63:0] X477;
   wire [63:0] Y477;
   wire [63:0] X478;
   wire [63:0] Y478;
   wire [63:0] X479;
   wire [63:0] Y479;
   wire [63:0] X480;
   wire [63:0] Y480;
   wire [63:0] X481;
   wire [63:0] Y481;
   wire [63:0] X482;
   wire [63:0] Y482;
   wire [63:0] X483;
   wire [63:0] Y483;
   wire [63:0] X484;
   wire [63:0] Y484;
   wire [63:0] X485;
   wire [63:0] Y485;
   wire [63:0] X486;
   wire [63:0] Y486;
   wire [63:0] X487;
   wire [63:0] Y487;
   wire [63:0] X488;
   wire [63:0] Y488;
   wire [63:0] X489;
   wire [63:0] Y489;
   wire [63:0] X490;
   wire [63:0] Y490;
   wire [63:0] X491;
   wire [63:0] Y491;
   wire [63:0] X492;
   wire [63:0] Y492;
   wire [63:0] X493;
   wire [63:0] Y493;
   wire [63:0] X494;
   wire [63:0] Y494;
   wire [63:0] X495;
   wire [63:0] Y495;
   wire [63:0] X496;
   wire [63:0] Y496;
   wire [63:0] X497;
   wire [63:0] Y497;
   wire [63:0] X498;
   wire [63:0] Y498;
   wire [63:0] X499;
   wire [63:0] Y499;
   wire [63:0] X500;
   wire [63:0] Y500;
   wire [63:0] X501;
   wire [63:0] Y501;
   wire [63:0] X502;
   wire [63:0] Y502;
   wire [63:0] X503;
   wire [63:0] Y503;
   wire [63:0] X504;
   wire [63:0] Y504;
   wire [63:0] X505;
   wire [63:0] Y505;
   wire [63:0] X506;
   wire [63:0] Y506;
   wire [63:0] X507;
   wire [63:0] Y507;
   wire [63:0] X508;
   wire [63:0] Y508;
   wire [63:0] X509;
   wire [63:0] Y509;
   wire [63:0] X510;
   wire [63:0] Y510;
   wire [63:0] X511;
   wire [63:0] Y511;
   wire [63:0] X512;
   wire [63:0] Y512;
   wire [63:0] X513;
   wire [63:0] Y513;
   wire [63:0] X514;
   wire [63:0] Y514;
   wire [63:0] X515;
   wire [63:0] Y515;
   wire [63:0] X516;
   wire [63:0] Y516;
   wire [63:0] X517;
   wire [63:0] Y517;
   wire [63:0] X518;
   wire [63:0] Y518;
   wire [63:0] X519;
   wire [63:0] Y519;
   wire [63:0] X520;
   wire [63:0] Y520;
   wire [63:0] X521;
   wire [63:0] Y521;
   wire [63:0] X522;
   wire [63:0] Y522;
   wire [63:0] X523;
   wire [63:0] Y523;
   wire [63:0] X524;
   wire [63:0] Y524;
   wire [63:0] X525;
   wire [63:0] Y525;
   wire [63:0] X526;
   wire [63:0] Y526;
   wire [63:0] X527;
   wire [63:0] Y527;
   wire [63:0] X528;
   wire [63:0] Y528;
   wire [63:0] X529;
   wire [63:0] Y529;
   wire [63:0] X530;
   wire [63:0] Y530;
   wire [63:0] X531;
   wire [63:0] Y531;
   wire [63:0] X532;
   wire [63:0] Y532;
   wire [63:0] X533;
   wire [63:0] Y533;
   wire [63:0] X534;
   wire [63:0] Y534;
   wire [63:0] X535;
   wire [63:0] Y535;
   wire [63:0] X536;
   wire [63:0] Y536;
   wire [63:0] X537;
   wire [63:0] Y537;
   wire [63:0] X538;
   wire [63:0] Y538;
   wire [63:0] X539;
   wire [63:0] Y539;
   wire [63:0] X540;
   wire [63:0] Y540;
   wire [63:0] X541;
   wire [63:0] Y541;
   wire [63:0] X542;
   wire [63:0] Y542;
   wire [63:0] X543;
   wire [63:0] Y543;
   wire [63:0] X544;
   wire [63:0] Y544;
   wire [63:0] X545;
   wire [63:0] Y545;
   wire [63:0] X546;
   wire [63:0] Y546;
   wire [63:0] X547;
   wire [63:0] Y547;
   wire [63:0] X548;
   wire [63:0] Y548;
   wire [63:0] X549;
   wire [63:0] Y549;
   wire [63:0] X550;
   wire [63:0] Y550;
   wire [63:0] X551;
   wire [63:0] Y551;
   wire [63:0] X552;
   wire [63:0] Y552;
   wire [63:0] X553;
   wire [63:0] Y553;
   wire [63:0] X554;
   wire [63:0] Y554;
   wire [63:0] X555;
   wire [63:0] Y555;
   wire [63:0] X556;
   wire [63:0] Y556;
   wire [63:0] X557;
   wire [63:0] Y557;
   wire [63:0] X558;
   wire [63:0] Y558;
   wire [63:0] X559;
   wire [63:0] Y559;
   wire [63:0] X560;
   wire [63:0] Y560;
   wire [63:0] X561;
   wire [63:0] Y561;
   wire [63:0] X562;
   wire [63:0] Y562;
   wire [63:0] X563;
   wire [63:0] Y563;
   wire [63:0] X564;
   wire [63:0] Y564;
   wire [63:0] X565;
   wire [63:0] Y565;
   wire [63:0] X566;
   wire [63:0] Y566;
   wire [63:0] X567;
   wire [63:0] Y567;
   wire [63:0] X568;
   wire [63:0] Y568;
   wire [63:0] X569;
   wire [63:0] Y569;
   wire [63:0] X570;
   wire [63:0] Y570;
   wire [63:0] X571;
   wire [63:0] Y571;
   wire [63:0] X572;
   wire [63:0] Y572;
   wire [63:0] X573;
   wire [63:0] Y573;
   wire [63:0] X574;
   wire [63:0] Y574;
   wire [63:0] X575;
   wire [63:0] Y575;
   wire [63:0] X576;
   wire [63:0] Y576;
   wire [63:0] X577;
   wire [63:0] Y577;
   wire [63:0] X578;
   wire [63:0] Y578;
   wire [63:0] X579;
   wire [63:0] Y579;
   wire [63:0] X580;
   wire [63:0] Y580;
   wire [63:0] X581;
   wire [63:0] Y581;
   wire [63:0] X582;
   wire [63:0] Y582;
   wire [63:0] X583;
   wire [63:0] Y583;
   wire [63:0] X584;
   wire [63:0] Y584;
   wire [63:0] X585;
   wire [63:0] Y585;
   wire [63:0] X586;
   wire [63:0] Y586;
   wire [63:0] X587;
   wire [63:0] Y587;
   wire [63:0] X588;
   wire [63:0] Y588;
   wire [63:0] X589;
   wire [63:0] Y589;
   wire [63:0] X590;
   wire [63:0] Y590;
   wire [63:0] X591;
   wire [63:0] Y591;
   wire [63:0] X592;
   wire [63:0] Y592;
   wire [63:0] X593;
   wire [63:0] Y593;
   wire [63:0] X594;
   wire [63:0] Y594;
   wire [63:0] X595;
   wire [63:0] Y595;
   wire [63:0] X596;
   wire [63:0] Y596;
   wire [63:0] X597;
   wire [63:0] Y597;
   wire [63:0] X598;
   wire [63:0] Y598;
   wire [63:0] X599;
   wire [63:0] Y599;
   wire [63:0] X600;
   wire [63:0] Y600;
   wire [63:0] X601;
   wire [63:0] Y601;
   wire [63:0] X602;
   wire [63:0] Y602;
   wire [63:0] X603;
   wire [63:0] Y603;
   wire [63:0] X604;
   wire [63:0] Y604;
   wire [63:0] X605;
   wire [63:0] Y605;
   wire [63:0] X606;
   wire [63:0] Y606;
   wire [63:0] X607;
   wire [63:0] Y607;
   wire [63:0] X608;
   wire [63:0] Y608;
   wire [63:0] X609;
   wire [63:0] Y609;
   wire [63:0] X610;
   wire [63:0] Y610;
   wire [63:0] X611;
   wire [63:0] Y611;
   wire [63:0] X612;
   wire [63:0] Y612;
   wire [63:0] X613;
   wire [63:0] Y613;
   wire [63:0] X614;
   wire [63:0] Y614;
   wire [63:0] X615;
   wire [63:0] Y615;
   wire [63:0] X616;
   wire [63:0] Y616;
   wire [63:0] X617;
   wire [63:0] Y617;
   wire [63:0] X618;
   wire [63:0] Y618;
   wire [63:0] X619;
   wire [63:0] Y619;
   wire [63:0] X620;
   wire [63:0] Y620;
   wire [63:0] X621;
   wire [63:0] Y621;
   wire [63:0] X622;
   wire [63:0] Y622;
   wire [63:0] X623;
   wire [63:0] Y623;
   wire [63:0] X624;
   wire [63:0] Y624;
   wire [63:0] X625;
   wire [63:0] Y625;
   wire [63:0] X626;
   wire [63:0] Y626;
   wire [63:0] X627;
   wire [63:0] Y627;
   wire [63:0] X628;
   wire [63:0] Y628;
   wire [63:0] X629;
   wire [63:0] Y629;
   wire [63:0] X630;
   wire [63:0] Y630;
   wire [63:0] X631;
   wire [63:0] Y631;
   wire [63:0] X632;
   wire [63:0] Y632;
   wire [63:0] X633;
   wire [63:0] Y633;
   wire [63:0] X634;
   wire [63:0] Y634;
   wire [63:0] X635;
   wire [63:0] Y635;
   wire [63:0] X636;
   wire [63:0] Y636;
   wire [63:0] X637;
   wire [63:0] Y637;
   wire [63:0] X638;
   wire [63:0] Y638;
   wire [63:0] X639;
   wire [63:0] Y639;
   wire [63:0] X640;
   wire [63:0] Y640;
   wire [63:0] X641;
   wire [63:0] Y641;
   wire [63:0] X642;
   wire [63:0] Y642;
   wire [63:0] X643;
   wire [63:0] Y643;
   wire [63:0] X644;
   wire [63:0] Y644;
   wire [63:0] X645;
   wire [63:0] Y645;
   wire [63:0] X646;
   wire [63:0] Y646;
   wire [63:0] X647;
   wire [63:0] Y647;
   wire [63:0] X648;
   wire [63:0] Y648;
   wire [63:0] X649;
   wire [63:0] Y649;
   wire [63:0] X650;
   wire [63:0] Y650;
   wire [63:0] X651;
   wire [63:0] Y651;
   wire [63:0] X652;
   wire [63:0] Y652;
   wire [63:0] X653;
   wire [63:0] Y653;
   wire [63:0] X654;
   wire [63:0] Y654;
   wire [63:0] X655;
   wire [63:0] Y655;
   wire [63:0] X656;
   wire [63:0] Y656;
   wire [63:0] X657;
   wire [63:0] Y657;
   wire [63:0] X658;
   wire [63:0] Y658;
   wire [63:0] X659;
   wire [63:0] Y659;
   wire [63:0] X660;
   wire [63:0] Y660;
   wire [63:0] X661;
   wire [63:0] Y661;
   wire [63:0] X662;
   wire [63:0] Y662;
   wire [63:0] X663;
   wire [63:0] Y663;
   wire [63:0] X664;
   wire [63:0] Y664;
   wire [63:0] X665;
   wire [63:0] Y665;
   wire [63:0] X666;
   wire [63:0] Y666;
   wire [63:0] X667;
   wire [63:0] Y667;
   wire [63:0] X668;
   wire [63:0] Y668;
   wire [63:0] X669;
   wire [63:0] Y669;
   wire [63:0] X670;
   wire [63:0] Y670;
   wire [63:0] X671;
   wire [63:0] Y671;
   wire [63:0] X672;
   wire [63:0] Y672;
   wire [63:0] X673;
   wire [63:0] Y673;
   wire [63:0] X674;
   wire [63:0] Y674;
   wire [63:0] X675;
   wire [63:0] Y675;
   wire [63:0] X676;
   wire [63:0] Y676;
   wire [63:0] X677;
   wire [63:0] Y677;
   wire [63:0] X678;
   wire [63:0] Y678;
   wire [63:0] X679;
   wire [63:0] Y679;
   wire [63:0] X680;
   wire [63:0] Y680;
   wire [63:0] X681;
   wire [63:0] Y681;
   wire [63:0] X682;
   wire [63:0] Y682;
   wire [63:0] X683;
   wire [63:0] Y683;
   wire [63:0] X684;
   wire [63:0] Y684;
   wire [63:0] X685;
   wire [63:0] Y685;
   wire [63:0] X686;
   wire [63:0] Y686;
   wire [63:0] X687;
   wire [63:0] Y687;
   wire [63:0] X688;
   wire [63:0] Y688;
   wire [63:0] X689;
   wire [63:0] Y689;
   wire [63:0] X690;
   wire [63:0] Y690;
   wire [63:0] X691;
   wire [63:0] Y691;
   wire [63:0] X692;
   wire [63:0] Y692;
   wire [63:0] X693;
   wire [63:0] Y693;
   wire [63:0] X694;
   wire [63:0] Y694;
   wire [63:0] X695;
   wire [63:0] Y695;
   wire [63:0] X696;
   wire [63:0] Y696;
   wire [63:0] X697;
   wire [63:0] Y697;
   wire [63:0] X698;
   wire [63:0] Y698;
   wire [63:0] X699;
   wire [63:0] Y699;
   wire [63:0] X700;
   wire [63:0] Y700;
   wire [63:0] X701;
   wire [63:0] Y701;
   wire [63:0] X702;
   wire [63:0] Y702;
   wire [63:0] X703;
   wire [63:0] Y703;
   wire [63:0] X704;
   wire [63:0] Y704;
   wire [63:0] X705;
   wire [63:0] Y705;
   wire [63:0] X706;
   wire [63:0] Y706;
   wire [63:0] X707;
   wire [63:0] Y707;
   wire [63:0] X708;
   wire [63:0] Y708;
   wire [63:0] X709;
   wire [63:0] Y709;
   wire [63:0] X710;
   wire [63:0] Y710;
   wire [63:0] X711;
   wire [63:0] Y711;
   wire [63:0] X712;
   wire [63:0] Y712;
   wire [63:0] X713;
   wire [63:0] Y713;
   wire [63:0] X714;
   wire [63:0] Y714;
   wire [63:0] X715;
   wire [63:0] Y715;
   wire [63:0] X716;
   wire [63:0] Y716;
   wire [63:0] X717;
   wire [63:0] Y717;
   wire [63:0] X718;
   wire [63:0] Y718;
   wire [63:0] X719;
   wire [63:0] Y719;
   wire [63:0] X720;
   wire [63:0] Y720;
   wire [63:0] X721;
   wire [63:0] Y721;
   wire [63:0] X722;
   wire [63:0] Y722;
   wire [63:0] X723;
   wire [63:0] Y723;
   wire [63:0] X724;
   wire [63:0] Y724;
   wire [63:0] X725;
   wire [63:0] Y725;
   wire [63:0] X726;
   wire [63:0] Y726;
   wire [63:0] X727;
   wire [63:0] Y727;
   wire [63:0] X728;
   wire [63:0] Y728;
   wire [63:0] X729;
   wire [63:0] Y729;
   wire [63:0] X730;
   wire [63:0] Y730;
   wire [63:0] X731;
   wire [63:0] Y731;
   wire [63:0] X732;
   wire [63:0] Y732;
   wire [63:0] X733;
   wire [63:0] Y733;
   wire [63:0] X734;
   wire [63:0] Y734;
   wire [63:0] X735;
   wire [63:0] Y735;
   wire [63:0] X736;
   wire [63:0] Y736;
   wire [63:0] X737;
   wire [63:0] Y737;
   wire [63:0] X738;
   wire [63:0] Y738;
   wire [63:0] X739;
   wire [63:0] Y739;
   wire [63:0] X740;
   wire [63:0] Y740;
   wire [63:0] X741;
   wire [63:0] Y741;
   wire [63:0] X742;
   wire [63:0] Y742;
   wire [63:0] X743;
   wire [63:0] Y743;
   wire [63:0] X744;
   wire [63:0] Y744;
   wire [63:0] X745;
   wire [63:0] Y745;
   wire [63:0] X746;
   wire [63:0] Y746;
   wire [63:0] X747;
   wire [63:0] Y747;
   wire [63:0] X748;
   wire [63:0] Y748;
   wire [63:0] X749;
   wire [63:0] Y749;
   wire [63:0] X750;
   wire [63:0] Y750;
   wire [63:0] X751;
   wire [63:0] Y751;
   wire [63:0] X752;
   wire [63:0] Y752;
   wire [63:0] X753;
   wire [63:0] Y753;
   wire [63:0] X754;
   wire [63:0] Y754;
   wire [63:0] X755;
   wire [63:0] Y755;
   wire [63:0] X756;
   wire [63:0] Y756;
   wire [63:0] X757;
   wire [63:0] Y757;
   wire [63:0] X758;
   wire [63:0] Y758;
   wire [63:0] X759;
   wire [63:0] Y759;
   wire [63:0] X760;
   wire [63:0] Y760;
   wire [63:0] X761;
   wire [63:0] Y761;
   wire [63:0] X762;
   wire [63:0] Y762;
   wire [63:0] X763;
   wire [63:0] Y763;
   wire [63:0] X764;
   wire [63:0] Y764;
   wire [63:0] X765;
   wire [63:0] Y765;
   wire [63:0] X766;
   wire [63:0] Y766;
   wire [63:0] X767;
   wire [63:0] Y767;
   wire [63:0] X768;
   wire [63:0] Y768;
   wire [63:0] X769;
   wire [63:0] Y769;
   wire [63:0] X770;
   wire [63:0] Y770;
   wire [63:0] X771;
   wire [63:0] Y771;
   wire [63:0] X772;
   wire [63:0] Y772;
   wire [63:0] X773;
   wire [63:0] Y773;
   wire [63:0] X774;
   wire [63:0] Y774;
   wire [63:0] X775;
   wire [63:0] Y775;
   wire [63:0] X776;
   wire [63:0] Y776;
   wire [63:0] X777;
   wire [63:0] Y777;
   wire [63:0] X778;
   wire [63:0] Y778;
   wire [63:0] X779;
   wire [63:0] Y779;
   wire [63:0] X780;
   wire [63:0] Y780;
   wire [63:0] X781;
   wire [63:0] Y781;
   wire [63:0] X782;
   wire [63:0] Y782;
   wire [63:0] X783;
   wire [63:0] Y783;
   wire [63:0] X784;
   wire [63:0] Y784;
   wire [63:0] X785;
   wire [63:0] Y785;
   wire [63:0] X786;
   wire [63:0] Y786;
   wire [63:0] X787;
   wire [63:0] Y787;
   wire [63:0] X788;
   wire [63:0] Y788;
   wire [63:0] X789;
   wire [63:0] Y789;
   wire [63:0] X790;
   wire [63:0] Y790;
   wire [63:0] X791;
   wire [63:0] Y791;
   wire [63:0] X792;
   wire [63:0] Y792;
   wire [63:0] X793;
   wire [63:0] Y793;
   wire [63:0] X794;
   wire [63:0] Y794;
   wire [63:0] X795;
   wire [63:0] Y795;
   wire [63:0] X796;
   wire [63:0] Y796;
   wire [63:0] X797;
   wire [63:0] Y797;
   wire [63:0] X798;
   wire [63:0] Y798;
   wire [63:0] X799;
   wire [63:0] Y799;
   wire [63:0] X800;
   wire [63:0] Y800;
   wire [63:0] X801;
   wire [63:0] Y801;
   wire [63:0] X802;
   wire [63:0] Y802;
   wire [63:0] X803;
   wire [63:0] Y803;
   wire [63:0] X804;
   wire [63:0] Y804;
   wire [63:0] X805;
   wire [63:0] Y805;
   wire [63:0] X806;
   wire [63:0] Y806;
   wire [63:0] X807;
   wire [63:0] Y807;
   wire [63:0] X808;
   wire [63:0] Y808;
   wire [63:0] X809;
   wire [63:0] Y809;
   wire [63:0] X810;
   wire [63:0] Y810;
   wire [63:0] X811;
   wire [63:0] Y811;
   wire [63:0] X812;
   wire [63:0] Y812;
   wire [63:0] X813;
   wire [63:0] Y813;
   wire [63:0] X814;
   wire [63:0] Y814;
   wire [63:0] X815;
   wire [63:0] Y815;
   wire [63:0] X816;
   wire [63:0] Y816;
   wire [63:0] X817;
   wire [63:0] Y817;
   wire [63:0] X818;
   wire [63:0] Y818;
   wire [63:0] X819;
   wire [63:0] Y819;
   wire [63:0] X820;
   wire [63:0] Y820;
   wire [63:0] X821;
   wire [63:0] Y821;
   wire [63:0] X822;
   wire [63:0] Y822;
   wire [63:0] X823;
   wire [63:0] Y823;
   wire [63:0] X824;
   wire [63:0] Y824;
   wire [63:0] X825;
   wire [63:0] Y825;
   wire [63:0] X826;
   wire [63:0] Y826;
   wire [63:0] X827;
   wire [63:0] Y827;
   wire [63:0] X828;
   wire [63:0] Y828;
   wire [63:0] X829;
   wire [63:0] Y829;
   wire [63:0] X830;
   wire [63:0] Y830;
   wire [63:0] X831;
   wire [63:0] Y831;
   wire [63:0] X832;
   wire [63:0] Y832;
   wire [63:0] X833;
   wire [63:0] Y833;
   wire [63:0] X834;
   wire [63:0] Y834;
   wire [63:0] X835;
   wire [63:0] Y835;
   wire [63:0] X836;
   wire [63:0] Y836;
   wire [63:0] X837;
   wire [63:0] Y837;
   wire [63:0] X838;
   wire [63:0] Y838;
   wire [63:0] X839;
   wire [63:0] Y839;
   wire [63:0] X840;
   wire [63:0] Y840;
   wire [63:0] X841;
   wire [63:0] Y841;
   wire [63:0] X842;
   wire [63:0] Y842;
   wire [63:0] X843;
   wire [63:0] Y843;
   wire [63:0] X844;
   wire [63:0] Y844;
   wire [63:0] X845;
   wire [63:0] Y845;
   wire [63:0] X846;
   wire [63:0] Y846;
   wire [63:0] X847;
   wire [63:0] Y847;
   wire [63:0] X848;
   wire [63:0] Y848;
   wire [63:0] X849;
   wire [63:0] Y849;
   wire [63:0] X850;
   wire [63:0] Y850;
   wire [63:0] X851;
   wire [63:0] Y851;
   wire [63:0] X852;
   wire [63:0] Y852;
   wire [63:0] X853;
   wire [63:0] Y853;
   wire [63:0] X854;
   wire [63:0] Y854;
   wire [63:0] X855;
   wire [63:0] Y855;
   wire [63:0] X856;
   wire [63:0] Y856;
   wire [63:0] X857;
   wire [63:0] Y857;
   wire [63:0] X858;
   wire [63:0] Y858;
   wire [63:0] X859;
   wire [63:0] Y859;
   wire [63:0] X860;
   wire [63:0] Y860;
   wire [63:0] X861;
   wire [63:0] Y861;
   wire [63:0] X862;
   wire [63:0] Y862;
   wire [63:0] X863;
   wire [63:0] Y863;
   wire [63:0] X864;
   wire [63:0] Y864;
   wire [63:0] X865;
   wire [63:0] Y865;
   wire [63:0] X866;
   wire [63:0] Y866;
   wire [63:0] X867;
   wire [63:0] Y867;
   wire [63:0] X868;
   wire [63:0] Y868;
   wire [63:0] X869;
   wire [63:0] Y869;
   wire [63:0] X870;
   wire [63:0] Y870;
   wire [63:0] X871;
   wire [63:0] Y871;
   wire [63:0] X872;
   wire [63:0] Y872;
   wire [63:0] X873;
   wire [63:0] Y873;
   wire [63:0] X874;
   wire [63:0] Y874;
   wire [63:0] X875;
   wire [63:0] Y875;
   wire [63:0] X876;
   wire [63:0] Y876;
   wire [63:0] X877;
   wire [63:0] Y877;
   wire [63:0] X878;
   wire [63:0] Y878;
   wire [63:0] X879;
   wire [63:0] Y879;
   wire [63:0] X880;
   wire [63:0] Y880;
   wire [63:0] X881;
   wire [63:0] Y881;
   wire [63:0] X882;
   wire [63:0] Y882;
   wire [63:0] X883;
   wire [63:0] Y883;
   wire [63:0] X884;
   wire [63:0] Y884;
   wire [63:0] X885;
   wire [63:0] Y885;
   wire [63:0] X886;
   wire [63:0] Y886;
   wire [63:0] X887;
   wire [63:0] Y887;
   wire [63:0] X888;
   wire [63:0] Y888;
   wire [63:0] X889;
   wire [63:0] Y889;
   wire [63:0] X890;
   wire [63:0] Y890;
   wire [63:0] X891;
   wire [63:0] Y891;
   wire [63:0] X892;
   wire [63:0] Y892;
   wire [63:0] X893;
   wire [63:0] Y893;
   wire [63:0] X894;
   wire [63:0] Y894;
   wire [63:0] X895;
   wire [63:0] Y895;
   wire [63:0] X896;
   wire [63:0] Y896;
   wire [63:0] X897;
   wire [63:0] Y897;
   wire [63:0] X898;
   wire [63:0] Y898;
   wire [63:0] X899;
   wire [63:0] Y899;
   wire [63:0] X900;
   wire [63:0] Y900;
   wire [63:0] X901;
   wire [63:0] Y901;
   wire [63:0] X902;
   wire [63:0] Y902;
   wire [63:0] X903;
   wire [63:0] Y903;
   wire [63:0] X904;
   wire [63:0] Y904;
   wire [63:0] X905;
   wire [63:0] Y905;
   wire [63:0] X906;
   wire [63:0] Y906;
   wire [63:0] X907;
   wire [63:0] Y907;
   wire [63:0] X908;
   wire [63:0] Y908;
   wire [63:0] X909;
   wire [63:0] Y909;
   wire [63:0] X910;
   wire [63:0] Y910;
   wire [63:0] X911;
   wire [63:0] Y911;
   wire [63:0] X912;
   wire [63:0] Y912;
   wire [63:0] X913;
   wire [63:0] Y913;
   wire [63:0] X914;
   wire [63:0] Y914;
   wire [63:0] X915;
   wire [63:0] Y915;
   wire [63:0] X916;
   wire [63:0] Y916;
   wire [63:0] X917;
   wire [63:0] Y917;
   wire [63:0] X918;
   wire [63:0] Y918;
   wire [63:0] X919;
   wire [63:0] Y919;
   wire [63:0] X920;
   wire [63:0] Y920;
   wire [63:0] X921;
   wire [63:0] Y921;
   wire [63:0] X922;
   wire [63:0] Y922;
   wire [63:0] X923;
   wire [63:0] Y923;
   wire [63:0] X924;
   wire [63:0] Y924;
   wire [63:0] X925;
   wire [63:0] Y925;
   wire [63:0] X926;
   wire [63:0] Y926;
   wire [63:0] X927;
   wire [63:0] Y927;
   wire [63:0] X928;
   wire [63:0] Y928;
   wire [63:0] X929;
   wire [63:0] Y929;
   wire [63:0] X930;
   wire [63:0] Y930;
   wire [63:0] X931;
   wire [63:0] Y931;
   wire [63:0] X932;
   wire [63:0] Y932;
   wire [63:0] X933;
   wire [63:0] Y933;
   wire [63:0] X934;
   wire [63:0] Y934;
   wire [63:0] X935;
   wire [63:0] Y935;
   wire [63:0] X936;
   wire [63:0] Y936;
   wire [63:0] X937;
   wire [63:0] Y937;
   wire [63:0] X938;
   wire [63:0] Y938;
   wire [63:0] X939;
   wire [63:0] Y939;
   wire [63:0] X940;
   wire [63:0] Y940;
   wire [63:0] X941;
   wire [63:0] Y941;
   wire [63:0] X942;
   wire [63:0] Y942;
   wire [63:0] X943;
   wire [63:0] Y943;
   wire [63:0] X944;
   wire [63:0] Y944;
   wire [63:0] X945;
   wire [63:0] Y945;
   wire [63:0] X946;
   wire [63:0] Y946;
   wire [63:0] X947;
   wire [63:0] Y947;
   wire [63:0] X948;
   wire [63:0] Y948;
   wire [63:0] X949;
   wire [63:0] Y949;
   wire [63:0] X950;
   wire [63:0] Y950;
   wire [63:0] X951;
   wire [63:0] Y951;
   wire [63:0] X952;
   wire [63:0] Y952;
   wire [63:0] X953;
   wire [63:0] Y953;
   wire [63:0] X954;
   wire [63:0] Y954;
   wire [63:0] X955;
   wire [63:0] Y955;
   wire [63:0] X956;
   wire [63:0] Y956;
   wire [63:0] X957;
   wire [63:0] Y957;
   wire [63:0] X958;
   wire [63:0] Y958;
   wire [63:0] X959;
   wire [63:0] Y959;
   wire [63:0] X960;
   wire [63:0] Y960;
   wire [63:0] X961;
   wire [63:0] Y961;
   wire [63:0] X962;
   wire [63:0] Y962;
   wire [63:0] X963;
   wire [63:0] Y963;
   wire [63:0] X964;
   wire [63:0] Y964;
   wire [63:0] X965;
   wire [63:0] Y965;
   wire [63:0] X966;
   wire [63:0] Y966;
   wire [63:0] X967;
   wire [63:0] Y967;
   wire [63:0] X968;
   wire [63:0] Y968;
   wire [63:0] X969;
   wire [63:0] Y969;
   wire [63:0] X970;
   wire [63:0] Y970;
   wire [63:0] X971;
   wire [63:0] Y971;
   wire [63:0] X972;
   wire [63:0] Y972;
   wire [63:0] X973;
   wire [63:0] Y973;
   wire [63:0] X974;
   wire [63:0] Y974;
   wire [63:0] X975;
   wire [63:0] Y975;
   wire [63:0] X976;
   wire [63:0] Y976;
   wire [63:0] X977;
   wire [63:0] Y977;
   wire [63:0] X978;
   wire [63:0] Y978;
   wire [63:0] X979;
   wire [63:0] Y979;
   wire [63:0] X980;
   wire [63:0] Y980;
   wire [63:0] X981;
   wire [63:0] Y981;
   wire [63:0] X982;
   wire [63:0] Y982;
   wire [63:0] X983;
   wire [63:0] Y983;
   wire [63:0] X984;
   wire [63:0] Y984;
   wire [63:0] X985;
   wire [63:0] Y985;
   wire [63:0] X986;
   wire [63:0] Y986;
   wire [63:0] X987;
   wire [63:0] Y987;
   wire [63:0] X988;
   wire [63:0] Y988;
   wire [63:0] X989;
   wire [63:0] Y989;
   wire [63:0] X990;
   wire [63:0] Y990;
   wire [63:0] X991;
   wire [63:0] Y991;
   wire [63:0] X992;
   wire [63:0] Y992;
   wire [63:0] X993;
   wire [63:0] Y993;
   wire [63:0] X994;
   wire [63:0] Y994;
   wire [63:0] X995;
   wire [63:0] Y995;
   wire [63:0] X996;
   wire [63:0] Y996;
   wire [63:0] X997;
   wire [63:0] Y997;
   wire [63:0] X998;
   wire [63:0] Y998;
   wire [63:0] X999;
   wire [63:0] Y999;
   wire [63:0] X1000;
   wire [63:0] Y1000;
   wire [63:0] X1001;
   wire [63:0] Y1001;
   wire [63:0] X1002;
   wire [63:0] Y1002;
   wire [63:0] X1003;
   wire [63:0] Y1003;
   wire [63:0] X1004;
   wire [63:0] Y1004;
   wire [63:0] X1005;
   wire [63:0] Y1005;
   wire [63:0] X1006;
   wire [63:0] Y1006;
   wire [63:0] X1007;
   wire [63:0] Y1007;
   wire [63:0] X1008;
   wire [63:0] Y1008;
   wire [63:0] X1009;
   wire [63:0] Y1009;
   wire [63:0] X1010;
   wire [63:0] Y1010;
   wire [63:0] X1011;
   wire [63:0] Y1011;
   wire [63:0] X1012;
   wire [63:0] Y1012;
   wire [63:0] X1013;
   wire [63:0] Y1013;
   wire [63:0] X1014;
   wire [63:0] Y1014;
   wire [63:0] X1015;
   wire [63:0] Y1015;
   wire [63:0] X1016;
   wire [63:0] Y1016;
   wire [63:0] X1017;
   wire [63:0] Y1017;
   wire [63:0] X1018;
   wire [63:0] Y1018;
   wire [63:0] X1019;
   wire [63:0] Y1019;
   wire [63:0] X1020;
   wire [63:0] Y1020;
   wire [63:0] X1021;
   wire [63:0] Y1021;
   wire [63:0] X1022;
   wire [63:0] Y1022;
   wire [63:0] X1023;
   wire [63:0] Y1023;
   reg clrCnt;
   assign X0 = in[0];
   assign X1 = in[1];
   assign X2 = in[2];
   assign X3 = in[3];
   assign X4 = in[4];
   assign X5 = in[5];
   assign X6 = in[6];
   assign X7 = in[7];
   assign X8 = in[8];
   assign X9 = in[9];
   assign X10 = in[10];
   assign X11 = in[11];
   assign X12 = in[12];
   assign X13 = in[13];
   assign X14 = in[14];
   assign X15 = in[15];
   assign X16 = in[16];
   assign X17 = in[17];
   assign X18 = in[18];
   assign X19 = in[19];
   assign X20 = in[20];
   assign X21 = in[21];
   assign X22 = in[22];
   assign X23 = in[23];
   assign X24 = in[24];
   assign X25 = in[25];
   assign X26 = in[26];
   assign X27 = in[27];
   assign X28 = in[28];
   assign X29 = in[29];
   assign X30 = in[30];
   assign X31 = in[31];
   assign X32 = in[32];
   assign X33 = in[33];
   assign X34 = in[34];
   assign X35 = in[35];
   assign X36 = in[36];
   assign X37 = in[37];
   assign X38 = in[38];
   assign X39 = in[39];
   assign X40 = in[40];
   assign X41 = in[41];
   assign X42 = in[42];
   assign X43 = in[43];
   assign X44 = in[44];
   assign X45 = in[45];
   assign X46 = in[46];
   assign X47 = in[47];
   assign X48 = in[48];
   assign X49 = in[49];
   assign X50 = in[50];
   assign X51 = in[51];
   assign X52 = in[52];
   assign X53 = in[53];
   assign X54 = in[54];
   assign X55 = in[55];
   assign X56 = in[56];
   assign X57 = in[57];
   assign X58 = in[58];
   assign X59 = in[59];
   assign X60 = in[60];
   assign X61 = in[61];
   assign X62 = in[62];
   assign X63 = in[63];
   assign X64 = in[64];
   assign X65 = in[65];
   assign X66 = in[66];
   assign X67 = in[67];
   assign X68 = in[68];
   assign X69 = in[69];
   assign X70 = in[70];
   assign X71 = in[71];
   assign X72 = in[72];
   assign X73 = in[73];
   assign X74 = in[74];
   assign X75 = in[75];
   assign X76 = in[76];
   assign X77 = in[77];
   assign X78 = in[78];
   assign X79 = in[79];
   assign X80 = in[80];
   assign X81 = in[81];
   assign X82 = in[82];
   assign X83 = in[83];
   assign X84 = in[84];
   assign X85 = in[85];
   assign X86 = in[86];
   assign X87 = in[87];
   assign X88 = in[88];
   assign X89 = in[89];
   assign X90 = in[90];
   assign X91 = in[91];
   assign X92 = in[92];
   assign X93 = in[93];
   assign X94 = in[94];
   assign X95 = in[95];
   assign X96 = in[96];
   assign X97 = in[97];
   assign X98 = in[98];
   assign X99 = in[99];
   assign X100 = in[100];
   assign X101 = in[101];
   assign X102 = in[102];
   assign X103 = in[103];
   assign X104 = in[104];
   assign X105 = in[105];
   assign X106 = in[106];
   assign X107 = in[107];
   assign X108 = in[108];
   assign X109 = in[109];
   assign X110 = in[110];
   assign X111 = in[111];
   assign X112 = in[112];
   assign X113 = in[113];
   assign X114 = in[114];
   assign X115 = in[115];
   assign X116 = in[116];
   assign X117 = in[117];
   assign X118 = in[118];
   assign X119 = in[119];
   assign X120 = in[120];
   assign X121 = in[121];
   assign X122 = in[122];
   assign X123 = in[123];
   assign X124 = in[124];
   assign X125 = in[125];
   assign X126 = in[126];
   assign X127 = in[127];
   assign X128 = in[128];
   assign X129 = in[129];
   assign X130 = in[130];
   assign X131 = in[131];
   assign X132 = in[132];
   assign X133 = in[133];
   assign X134 = in[134];
   assign X135 = in[135];
   assign X136 = in[136];
   assign X137 = in[137];
   assign X138 = in[138];
   assign X139 = in[139];
   assign X140 = in[140];
   assign X141 = in[141];
   assign X142 = in[142];
   assign X143 = in[143];
   assign X144 = in[144];
   assign X145 = in[145];
   assign X146 = in[146];
   assign X147 = in[147];
   assign X148 = in[148];
   assign X149 = in[149];
   assign X150 = in[150];
   assign X151 = in[151];
   assign X152 = in[152];
   assign X153 = in[153];
   assign X154 = in[154];
   assign X155 = in[155];
   assign X156 = in[156];
   assign X157 = in[157];
   assign X158 = in[158];
   assign X159 = in[159];
   assign X160 = in[160];
   assign X161 = in[161];
   assign X162 = in[162];
   assign X163 = in[163];
   assign X164 = in[164];
   assign X165 = in[165];
   assign X166 = in[166];
   assign X167 = in[167];
   assign X168 = in[168];
   assign X169 = in[169];
   assign X170 = in[170];
   assign X171 = in[171];
   assign X172 = in[172];
   assign X173 = in[173];
   assign X174 = in[174];
   assign X175 = in[175];
   assign X176 = in[176];
   assign X177 = in[177];
   assign X178 = in[178];
   assign X179 = in[179];
   assign X180 = in[180];
   assign X181 = in[181];
   assign X182 = in[182];
   assign X183 = in[183];
   assign X184 = in[184];
   assign X185 = in[185];
   assign X186 = in[186];
   assign X187 = in[187];
   assign X188 = in[188];
   assign X189 = in[189];
   assign X190 = in[190];
   assign X191 = in[191];
   assign X192 = in[192];
   assign X193 = in[193];
   assign X194 = in[194];
   assign X195 = in[195];
   assign X196 = in[196];
   assign X197 = in[197];
   assign X198 = in[198];
   assign X199 = in[199];
   assign X200 = in[200];
   assign X201 = in[201];
   assign X202 = in[202];
   assign X203 = in[203];
   assign X204 = in[204];
   assign X205 = in[205];
   assign X206 = in[206];
   assign X207 = in[207];
   assign X208 = in[208];
   assign X209 = in[209];
   assign X210 = in[210];
   assign X211 = in[211];
   assign X212 = in[212];
   assign X213 = in[213];
   assign X214 = in[214];
   assign X215 = in[215];
   assign X216 = in[216];
   assign X217 = in[217];
   assign X218 = in[218];
   assign X219 = in[219];
   assign X220 = in[220];
   assign X221 = in[221];
   assign X222 = in[222];
   assign X223 = in[223];
   assign X224 = in[224];
   assign X225 = in[225];
   assign X226 = in[226];
   assign X227 = in[227];
   assign X228 = in[228];
   assign X229 = in[229];
   assign X230 = in[230];
   assign X231 = in[231];
   assign X232 = in[232];
   assign X233 = in[233];
   assign X234 = in[234];
   assign X235 = in[235];
   assign X236 = in[236];
   assign X237 = in[237];
   assign X238 = in[238];
   assign X239 = in[239];
   assign X240 = in[240];
   assign X241 = in[241];
   assign X242 = in[242];
   assign X243 = in[243];
   assign X244 = in[244];
   assign X245 = in[245];
   assign X246 = in[246];
   assign X247 = in[247];
   assign X248 = in[248];
   assign X249 = in[249];
   assign X250 = in[250];
   assign X251 = in[251];
   assign X252 = in[252];
   assign X253 = in[253];
   assign X254 = in[254];
   assign X255 = in[255];
   assign X256 = in[256];
   assign X257 = in[257];
   assign X258 = in[258];
   assign X259 = in[259];
   assign X260 = in[260];
   assign X261 = in[261];
   assign X262 = in[262];
   assign X263 = in[263];
   assign X264 = in[264];
   assign X265 = in[265];
   assign X266 = in[266];
   assign X267 = in[267];
   assign X268 = in[268];
   assign X269 = in[269];
   assign X270 = in[270];
   assign X271 = in[271];
   assign X272 = in[272];
   assign X273 = in[273];
   assign X274 = in[274];
   assign X275 = in[275];
   assign X276 = in[276];
   assign X277 = in[277];
   assign X278 = in[278];
   assign X279 = in[279];
   assign X280 = in[280];
   assign X281 = in[281];
   assign X282 = in[282];
   assign X283 = in[283];
   assign X284 = in[284];
   assign X285 = in[285];
   assign X286 = in[286];
   assign X287 = in[287];
   assign X288 = in[288];
   assign X289 = in[289];
   assign X290 = in[290];
   assign X291 = in[291];
   assign X292 = in[292];
   assign X293 = in[293];
   assign X294 = in[294];
   assign X295 = in[295];
   assign X296 = in[296];
   assign X297 = in[297];
   assign X298 = in[298];
   assign X299 = in[299];
   assign X300 = in[300];
   assign X301 = in[301];
   assign X302 = in[302];
   assign X303 = in[303];
   assign X304 = in[304];
   assign X305 = in[305];
   assign X306 = in[306];
   assign X307 = in[307];
   assign X308 = in[308];
   assign X309 = in[309];
   assign X310 = in[310];
   assign X311 = in[311];
   assign X312 = in[312];
   assign X313 = in[313];
   assign X314 = in[314];
   assign X315 = in[315];
   assign X316 = in[316];
   assign X317 = in[317];
   assign X318 = in[318];
   assign X319 = in[319];
   assign X320 = in[320];
   assign X321 = in[321];
   assign X322 = in[322];
   assign X323 = in[323];
   assign X324 = in[324];
   assign X325 = in[325];
   assign X326 = in[326];
   assign X327 = in[327];
   assign X328 = in[328];
   assign X329 = in[329];
   assign X330 = in[330];
   assign X331 = in[331];
   assign X332 = in[332];
   assign X333 = in[333];
   assign X334 = in[334];
   assign X335 = in[335];
   assign X336 = in[336];
   assign X337 = in[337];
   assign X338 = in[338];
   assign X339 = in[339];
   assign X340 = in[340];
   assign X341 = in[341];
   assign X342 = in[342];
   assign X343 = in[343];
   assign X344 = in[344];
   assign X345 = in[345];
   assign X346 = in[346];
   assign X347 = in[347];
   assign X348 = in[348];
   assign X349 = in[349];
   assign X350 = in[350];
   assign X351 = in[351];
   assign X352 = in[352];
   assign X353 = in[353];
   assign X354 = in[354];
   assign X355 = in[355];
   assign X356 = in[356];
   assign X357 = in[357];
   assign X358 = in[358];
   assign X359 = in[359];
   assign X360 = in[360];
   assign X361 = in[361];
   assign X362 = in[362];
   assign X363 = in[363];
   assign X364 = in[364];
   assign X365 = in[365];
   assign X366 = in[366];
   assign X367 = in[367];
   assign X368 = in[368];
   assign X369 = in[369];
   assign X370 = in[370];
   assign X371 = in[371];
   assign X372 = in[372];
   assign X373 = in[373];
   assign X374 = in[374];
   assign X375 = in[375];
   assign X376 = in[376];
   assign X377 = in[377];
   assign X378 = in[378];
   assign X379 = in[379];
   assign X380 = in[380];
   assign X381 = in[381];
   assign X382 = in[382];
   assign X383 = in[383];
   assign X384 = in[384];
   assign X385 = in[385];
   assign X386 = in[386];
   assign X387 = in[387];
   assign X388 = in[388];
   assign X389 = in[389];
   assign X390 = in[390];
   assign X391 = in[391];
   assign X392 = in[392];
   assign X393 = in[393];
   assign X394 = in[394];
   assign X395 = in[395];
   assign X396 = in[396];
   assign X397 = in[397];
   assign X398 = in[398];
   assign X399 = in[399];
   assign X400 = in[400];
   assign X401 = in[401];
   assign X402 = in[402];
   assign X403 = in[403];
   assign X404 = in[404];
   assign X405 = in[405];
   assign X406 = in[406];
   assign X407 = in[407];
   assign X408 = in[408];
   assign X409 = in[409];
   assign X410 = in[410];
   assign X411 = in[411];
   assign X412 = in[412];
   assign X413 = in[413];
   assign X414 = in[414];
   assign X415 = in[415];
   assign X416 = in[416];
   assign X417 = in[417];
   assign X418 = in[418];
   assign X419 = in[419];
   assign X420 = in[420];
   assign X421 = in[421];
   assign X422 = in[422];
   assign X423 = in[423];
   assign X424 = in[424];
   assign X425 = in[425];
   assign X426 = in[426];
   assign X427 = in[427];
   assign X428 = in[428];
   assign X429 = in[429];
   assign X430 = in[430];
   assign X431 = in[431];
   assign X432 = in[432];
   assign X433 = in[433];
   assign X434 = in[434];
   assign X435 = in[435];
   assign X436 = in[436];
   assign X437 = in[437];
   assign X438 = in[438];
   assign X439 = in[439];
   assign X440 = in[440];
   assign X441 = in[441];
   assign X442 = in[442];
   assign X443 = in[443];
   assign X444 = in[444];
   assign X445 = in[445];
   assign X446 = in[446];
   assign X447 = in[447];
   assign X448 = in[448];
   assign X449 = in[449];
   assign X450 = in[450];
   assign X451 = in[451];
   assign X452 = in[452];
   assign X453 = in[453];
   assign X454 = in[454];
   assign X455 = in[455];
   assign X456 = in[456];
   assign X457 = in[457];
   assign X458 = in[458];
   assign X459 = in[459];
   assign X460 = in[460];
   assign X461 = in[461];
   assign X462 = in[462];
   assign X463 = in[463];
   assign X464 = in[464];
   assign X465 = in[465];
   assign X466 = in[466];
   assign X467 = in[467];
   assign X468 = in[468];
   assign X469 = in[469];
   assign X470 = in[470];
   assign X471 = in[471];
   assign X472 = in[472];
   assign X473 = in[473];
   assign X474 = in[474];
   assign X475 = in[475];
   assign X476 = in[476];
   assign X477 = in[477];
   assign X478 = in[478];
   assign X479 = in[479];
   assign X480 = in[480];
   assign X481 = in[481];
   assign X482 = in[482];
   assign X483 = in[483];
   assign X484 = in[484];
   assign X485 = in[485];
   assign X486 = in[486];
   assign X487 = in[487];
   assign X488 = in[488];
   assign X489 = in[489];
   assign X490 = in[490];
   assign X491 = in[491];
   assign X492 = in[492];
   assign X493 = in[493];
   assign X494 = in[494];
   assign X495 = in[495];
   assign X496 = in[496];
   assign X497 = in[497];
   assign X498 = in[498];
   assign X499 = in[499];
   assign X500 = in[500];
   assign X501 = in[501];
   assign X502 = in[502];
   assign X503 = in[503];
   assign X504 = in[504];
   assign X505 = in[505];
   assign X506 = in[506];
   assign X507 = in[507];
   assign X508 = in[508];
   assign X509 = in[509];
   assign X510 = in[510];
   assign X511 = in[511];
   assign X512 = in[512];
   assign X513 = in[513];
   assign X514 = in[514];
   assign X515 = in[515];
   assign X516 = in[516];
   assign X517 = in[517];
   assign X518 = in[518];
   assign X519 = in[519];
   assign X520 = in[520];
   assign X521 = in[521];
   assign X522 = in[522];
   assign X523 = in[523];
   assign X524 = in[524];
   assign X525 = in[525];
   assign X526 = in[526];
   assign X527 = in[527];
   assign X528 = in[528];
   assign X529 = in[529];
   assign X530 = in[530];
   assign X531 = in[531];
   assign X532 = in[532];
   assign X533 = in[533];
   assign X534 = in[534];
   assign X535 = in[535];
   assign X536 = in[536];
   assign X537 = in[537];
   assign X538 = in[538];
   assign X539 = in[539];
   assign X540 = in[540];
   assign X541 = in[541];
   assign X542 = in[542];
   assign X543 = in[543];
   assign X544 = in[544];
   assign X545 = in[545];
   assign X546 = in[546];
   assign X547 = in[547];
   assign X548 = in[548];
   assign X549 = in[549];
   assign X550 = in[550];
   assign X551 = in[551];
   assign X552 = in[552];
   assign X553 = in[553];
   assign X554 = in[554];
   assign X555 = in[555];
   assign X556 = in[556];
   assign X557 = in[557];
   assign X558 = in[558];
   assign X559 = in[559];
   assign X560 = in[560];
   assign X561 = in[561];
   assign X562 = in[562];
   assign X563 = in[563];
   assign X564 = in[564];
   assign X565 = in[565];
   assign X566 = in[566];
   assign X567 = in[567];
   assign X568 = in[568];
   assign X569 = in[569];
   assign X570 = in[570];
   assign X571 = in[571];
   assign X572 = in[572];
   assign X573 = in[573];
   assign X574 = in[574];
   assign X575 = in[575];
   assign X576 = in[576];
   assign X577 = in[577];
   assign X578 = in[578];
   assign X579 = in[579];
   assign X580 = in[580];
   assign X581 = in[581];
   assign X582 = in[582];
   assign X583 = in[583];
   assign X584 = in[584];
   assign X585 = in[585];
   assign X586 = in[586];
   assign X587 = in[587];
   assign X588 = in[588];
   assign X589 = in[589];
   assign X590 = in[590];
   assign X591 = in[591];
   assign X592 = in[592];
   assign X593 = in[593];
   assign X594 = in[594];
   assign X595 = in[595];
   assign X596 = in[596];
   assign X597 = in[597];
   assign X598 = in[598];
   assign X599 = in[599];
   assign X600 = in[600];
   assign X601 = in[601];
   assign X602 = in[602];
   assign X603 = in[603];
   assign X604 = in[604];
   assign X605 = in[605];
   assign X606 = in[606];
   assign X607 = in[607];
   assign X608 = in[608];
   assign X609 = in[609];
   assign X610 = in[610];
   assign X611 = in[611];
   assign X612 = in[612];
   assign X613 = in[613];
   assign X614 = in[614];
   assign X615 = in[615];
   assign X616 = in[616];
   assign X617 = in[617];
   assign X618 = in[618];
   assign X619 = in[619];
   assign X620 = in[620];
   assign X621 = in[621];
   assign X622 = in[622];
   assign X623 = in[623];
   assign X624 = in[624];
   assign X625 = in[625];
   assign X626 = in[626];
   assign X627 = in[627];
   assign X628 = in[628];
   assign X629 = in[629];
   assign X630 = in[630];
   assign X631 = in[631];
   assign X632 = in[632];
   assign X633 = in[633];
   assign X634 = in[634];
   assign X635 = in[635];
   assign X636 = in[636];
   assign X637 = in[637];
   assign X638 = in[638];
   assign X639 = in[639];
   assign X640 = in[640];
   assign X641 = in[641];
   assign X642 = in[642];
   assign X643 = in[643];
   assign X644 = in[644];
   assign X645 = in[645];
   assign X646 = in[646];
   assign X647 = in[647];
   assign X648 = in[648];
   assign X649 = in[649];
   assign X650 = in[650];
   assign X651 = in[651];
   assign X652 = in[652];
   assign X653 = in[653];
   assign X654 = in[654];
   assign X655 = in[655];
   assign X656 = in[656];
   assign X657 = in[657];
   assign X658 = in[658];
   assign X659 = in[659];
   assign X660 = in[660];
   assign X661 = in[661];
   assign X662 = in[662];
   assign X663 = in[663];
   assign X664 = in[664];
   assign X665 = in[665];
   assign X666 = in[666];
   assign X667 = in[667];
   assign X668 = in[668];
   assign X669 = in[669];
   assign X670 = in[670];
   assign X671 = in[671];
   assign X672 = in[672];
   assign X673 = in[673];
   assign X674 = in[674];
   assign X675 = in[675];
   assign X676 = in[676];
   assign X677 = in[677];
   assign X678 = in[678];
   assign X679 = in[679];
   assign X680 = in[680];
   assign X681 = in[681];
   assign X682 = in[682];
   assign X683 = in[683];
   assign X684 = in[684];
   assign X685 = in[685];
   assign X686 = in[686];
   assign X687 = in[687];
   assign X688 = in[688];
   assign X689 = in[689];
   assign X690 = in[690];
   assign X691 = in[691];
   assign X692 = in[692];
   assign X693 = in[693];
   assign X694 = in[694];
   assign X695 = in[695];
   assign X696 = in[696];
   assign X697 = in[697];
   assign X698 = in[698];
   assign X699 = in[699];
   assign X700 = in[700];
   assign X701 = in[701];
   assign X702 = in[702];
   assign X703 = in[703];
   assign X704 = in[704];
   assign X705 = in[705];
   assign X706 = in[706];
   assign X707 = in[707];
   assign X708 = in[708];
   assign X709 = in[709];
   assign X710 = in[710];
   assign X711 = in[711];
   assign X712 = in[712];
   assign X713 = in[713];
   assign X714 = in[714];
   assign X715 = in[715];
   assign X716 = in[716];
   assign X717 = in[717];
   assign X718 = in[718];
   assign X719 = in[719];
   assign X720 = in[720];
   assign X721 = in[721];
   assign X722 = in[722];
   assign X723 = in[723];
   assign X724 = in[724];
   assign X725 = in[725];
   assign X726 = in[726];
   assign X727 = in[727];
   assign X728 = in[728];
   assign X729 = in[729];
   assign X730 = in[730];
   assign X731 = in[731];
   assign X732 = in[732];
   assign X733 = in[733];
   assign X734 = in[734];
   assign X735 = in[735];
   assign X736 = in[736];
   assign X737 = in[737];
   assign X738 = in[738];
   assign X739 = in[739];
   assign X740 = in[740];
   assign X741 = in[741];
   assign X742 = in[742];
   assign X743 = in[743];
   assign X744 = in[744];
   assign X745 = in[745];
   assign X746 = in[746];
   assign X747 = in[747];
   assign X748 = in[748];
   assign X749 = in[749];
   assign X750 = in[750];
   assign X751 = in[751];
   assign X752 = in[752];
   assign X753 = in[753];
   assign X754 = in[754];
   assign X755 = in[755];
   assign X756 = in[756];
   assign X757 = in[757];
   assign X758 = in[758];
   assign X759 = in[759];
   assign X760 = in[760];
   assign X761 = in[761];
   assign X762 = in[762];
   assign X763 = in[763];
   assign X764 = in[764];
   assign X765 = in[765];
   assign X766 = in[766];
   assign X767 = in[767];
   assign X768 = in[768];
   assign X769 = in[769];
   assign X770 = in[770];
   assign X771 = in[771];
   assign X772 = in[772];
   assign X773 = in[773];
   assign X774 = in[774];
   assign X775 = in[775];
   assign X776 = in[776];
   assign X777 = in[777];
   assign X778 = in[778];
   assign X779 = in[779];
   assign X780 = in[780];
   assign X781 = in[781];
   assign X782 = in[782];
   assign X783 = in[783];
   assign X784 = in[784];
   assign X785 = in[785];
   assign X786 = in[786];
   assign X787 = in[787];
   assign X788 = in[788];
   assign X789 = in[789];
   assign X790 = in[790];
   assign X791 = in[791];
   assign X792 = in[792];
   assign X793 = in[793];
   assign X794 = in[794];
   assign X795 = in[795];
   assign X796 = in[796];
   assign X797 = in[797];
   assign X798 = in[798];
   assign X799 = in[799];
   assign X800 = in[800];
   assign X801 = in[801];
   assign X802 = in[802];
   assign X803 = in[803];
   assign X804 = in[804];
   assign X805 = in[805];
   assign X806 = in[806];
   assign X807 = in[807];
   assign X808 = in[808];
   assign X809 = in[809];
   assign X810 = in[810];
   assign X811 = in[811];
   assign X812 = in[812];
   assign X813 = in[813];
   assign X814 = in[814];
   assign X815 = in[815];
   assign X816 = in[816];
   assign X817 = in[817];
   assign X818 = in[818];
   assign X819 = in[819];
   assign X820 = in[820];
   assign X821 = in[821];
   assign X822 = in[822];
   assign X823 = in[823];
   assign X824 = in[824];
   assign X825 = in[825];
   assign X826 = in[826];
   assign X827 = in[827];
   assign X828 = in[828];
   assign X829 = in[829];
   assign X830 = in[830];
   assign X831 = in[831];
   assign X832 = in[832];
   assign X833 = in[833];
   assign X834 = in[834];
   assign X835 = in[835];
   assign X836 = in[836];
   assign X837 = in[837];
   assign X838 = in[838];
   assign X839 = in[839];
   assign X840 = in[840];
   assign X841 = in[841];
   assign X842 = in[842];
   assign X843 = in[843];
   assign X844 = in[844];
   assign X845 = in[845];
   assign X846 = in[846];
   assign X847 = in[847];
   assign X848 = in[848];
   assign X849 = in[849];
   assign X850 = in[850];
   assign X851 = in[851];
   assign X852 = in[852];
   assign X853 = in[853];
   assign X854 = in[854];
   assign X855 = in[855];
   assign X856 = in[856];
   assign X857 = in[857];
   assign X858 = in[858];
   assign X859 = in[859];
   assign X860 = in[860];
   assign X861 = in[861];
   assign X862 = in[862];
   assign X863 = in[863];
   assign X864 = in[864];
   assign X865 = in[865];
   assign X866 = in[866];
   assign X867 = in[867];
   assign X868 = in[868];
   assign X869 = in[869];
   assign X870 = in[870];
   assign X871 = in[871];
   assign X872 = in[872];
   assign X873 = in[873];
   assign X874 = in[874];
   assign X875 = in[875];
   assign X876 = in[876];
   assign X877 = in[877];
   assign X878 = in[878];
   assign X879 = in[879];
   assign X880 = in[880];
   assign X881 = in[881];
   assign X882 = in[882];
   assign X883 = in[883];
   assign X884 = in[884];
   assign X885 = in[885];
   assign X886 = in[886];
   assign X887 = in[887];
   assign X888 = in[888];
   assign X889 = in[889];
   assign X890 = in[890];
   assign X891 = in[891];
   assign X892 = in[892];
   assign X893 = in[893];
   assign X894 = in[894];
   assign X895 = in[895];
   assign X896 = in[896];
   assign X897 = in[897];
   assign X898 = in[898];
   assign X899 = in[899];
   assign X900 = in[900];
   assign X901 = in[901];
   assign X902 = in[902];
   assign X903 = in[903];
   assign X904 = in[904];
   assign X905 = in[905];
   assign X906 = in[906];
   assign X907 = in[907];
   assign X908 = in[908];
   assign X909 = in[909];
   assign X910 = in[910];
   assign X911 = in[911];
   assign X912 = in[912];
   assign X913 = in[913];
   assign X914 = in[914];
   assign X915 = in[915];
   assign X916 = in[916];
   assign X917 = in[917];
   assign X918 = in[918];
   assign X919 = in[919];
   assign X920 = in[920];
   assign X921 = in[921];
   assign X922 = in[922];
   assign X923 = in[923];
   assign X924 = in[924];
   assign X925 = in[925];
   assign X926 = in[926];
   assign X927 = in[927];
   assign X928 = in[928];
   assign X929 = in[929];
   assign X930 = in[930];
   assign X931 = in[931];
   assign X932 = in[932];
   assign X933 = in[933];
   assign X934 = in[934];
   assign X935 = in[935];
   assign X936 = in[936];
   assign X937 = in[937];
   assign X938 = in[938];
   assign X939 = in[939];
   assign X940 = in[940];
   assign X941 = in[941];
   assign X942 = in[942];
   assign X943 = in[943];
   assign X944 = in[944];
   assign X945 = in[945];
   assign X946 = in[946];
   assign X947 = in[947];
   assign X948 = in[948];
   assign X949 = in[949];
   assign X950 = in[950];
   assign X951 = in[951];
   assign X952 = in[952];
   assign X953 = in[953];
   assign X954 = in[954];
   assign X955 = in[955];
   assign X956 = in[956];
   assign X957 = in[957];
   assign X958 = in[958];
   assign X959 = in[959];
   assign X960 = in[960];
   assign X961 = in[961];
   assign X962 = in[962];
   assign X963 = in[963];
   assign X964 = in[964];
   assign X965 = in[965];
   assign X966 = in[966];
   assign X967 = in[967];
   assign X968 = in[968];
   assign X969 = in[969];
   assign X970 = in[970];
   assign X971 = in[971];
   assign X972 = in[972];
   assign X973 = in[973];
   assign X974 = in[974];
   assign X975 = in[975];
   assign X976 = in[976];
   assign X977 = in[977];
   assign X978 = in[978];
   assign X979 = in[979];
   assign X980 = in[980];
   assign X981 = in[981];
   assign X982 = in[982];
   assign X983 = in[983];
   assign X984 = in[984];
   assign X985 = in[985];
   assign X986 = in[986];
   assign X987 = in[987];
   assign X988 = in[988];
   assign X989 = in[989];
   assign X990 = in[990];
   assign X991 = in[991];
   assign X992 = in[992];
   assign X993 = in[993];
   assign X994 = in[994];
   assign X995 = in[995];
   assign X996 = in[996];
   assign X997 = in[997];
   assign X998 = in[998];
   assign X999 = in[999];
   assign X1000 = in[1000];
   assign X1001 = in[1001];
   assign X1002 = in[1002];
   assign X1003 = in[1003];
   assign X1004 = in[1004];
   assign X1005 = in[1005];
   assign X1006 = in[1006];
   assign X1007 = in[1007];
   assign X1008 = in[1008];
   assign X1009 = in[1009];
   assign X1010 = in[1010];
   assign X1011 = in[1011];
   assign X1012 = in[1012];
   assign X1013 = in[1013];
   assign X1014 = in[1014];
   assign X1015 = in[1015];
   assign X1016 = in[1016];
   assign X1017 = in[1017];
   assign X1018 = in[1018];
   assign X1019 = in[1019];
   assign X1020 = in[1020];
   assign X1021 = in[1021];
   assign X1022 = in[1022];
   assign X1023 = in[1023];

   initial clk = 0;

   always #10000 clk = ~clk;


   // Instantiate top-level module of core 'X' signals are system inputs
   // and 'Y' signals are system outputs
   dft_top dft_top_instance (.clk(clk), .reset(reset), .next(next), .next_out(next_out),
    .X0(X0), .Y0(Y0),
    .X1(X1), .Y1(Y1),
    .X2(X2), .Y2(Y2),
    .X3(X3), .Y3(Y3),
    .X4(X4), .Y4(Y4),
    .X5(X5), .Y5(Y5),
    .X6(X6), .Y6(Y6),
    .X7(X7), .Y7(Y7),
    .X8(X8), .Y8(Y8),
    .X9(X9), .Y9(Y9),
    .X10(X10), .Y10(Y10),
    .X11(X11), .Y11(Y11),
    .X12(X12), .Y12(Y12),
    .X13(X13), .Y13(Y13),
    .X14(X14), .Y14(Y14),
    .X15(X15), .Y15(Y15),
    .X16(X16), .Y16(Y16),
    .X17(X17), .Y17(Y17),
    .X18(X18), .Y18(Y18),
    .X19(X19), .Y19(Y19),
    .X20(X20), .Y20(Y20),
    .X21(X21), .Y21(Y21),
    .X22(X22), .Y22(Y22),
    .X23(X23), .Y23(Y23),
    .X24(X24), .Y24(Y24),
    .X25(X25), .Y25(Y25),
    .X26(X26), .Y26(Y26),
    .X27(X27), .Y27(Y27),
    .X28(X28), .Y28(Y28),
    .X29(X29), .Y29(Y29),
    .X30(X30), .Y30(Y30),
    .X31(X31), .Y31(Y31),
    .X32(X32), .Y32(Y32),
    .X33(X33), .Y33(Y33),
    .X34(X34), .Y34(Y34),
    .X35(X35), .Y35(Y35),
    .X36(X36), .Y36(Y36),
    .X37(X37), .Y37(Y37),
    .X38(X38), .Y38(Y38),
    .X39(X39), .Y39(Y39),
    .X40(X40), .Y40(Y40),
    .X41(X41), .Y41(Y41),
    .X42(X42), .Y42(Y42),
    .X43(X43), .Y43(Y43),
    .X44(X44), .Y44(Y44),
    .X45(X45), .Y45(Y45),
    .X46(X46), .Y46(Y46),
    .X47(X47), .Y47(Y47),
    .X48(X48), .Y48(Y48),
    .X49(X49), .Y49(Y49),
    .X50(X50), .Y50(Y50),
    .X51(X51), .Y51(Y51),
    .X52(X52), .Y52(Y52),
    .X53(X53), .Y53(Y53),
    .X54(X54), .Y54(Y54),
    .X55(X55), .Y55(Y55),
    .X56(X56), .Y56(Y56),
    .X57(X57), .Y57(Y57),
    .X58(X58), .Y58(Y58),
    .X59(X59), .Y59(Y59),
    .X60(X60), .Y60(Y60),
    .X61(X61), .Y61(Y61),
    .X62(X62), .Y62(Y62),
    .X63(X63), .Y63(Y63),
    .X64(X64), .Y64(Y64),
    .X65(X65), .Y65(Y65),
    .X66(X66), .Y66(Y66),
    .X67(X67), .Y67(Y67),
    .X68(X68), .Y68(Y68),
    .X69(X69), .Y69(Y69),
    .X70(X70), .Y70(Y70),
    .X71(X71), .Y71(Y71),
    .X72(X72), .Y72(Y72),
    .X73(X73), .Y73(Y73),
    .X74(X74), .Y74(Y74),
    .X75(X75), .Y75(Y75),
    .X76(X76), .Y76(Y76),
    .X77(X77), .Y77(Y77),
    .X78(X78), .Y78(Y78),
    .X79(X79), .Y79(Y79),
    .X80(X80), .Y80(Y80),
    .X81(X81), .Y81(Y81),
    .X82(X82), .Y82(Y82),
    .X83(X83), .Y83(Y83),
    .X84(X84), .Y84(Y84),
    .X85(X85), .Y85(Y85),
    .X86(X86), .Y86(Y86),
    .X87(X87), .Y87(Y87),
    .X88(X88), .Y88(Y88),
    .X89(X89), .Y89(Y89),
    .X90(X90), .Y90(Y90),
    .X91(X91), .Y91(Y91),
    .X92(X92), .Y92(Y92),
    .X93(X93), .Y93(Y93),
    .X94(X94), .Y94(Y94),
    .X95(X95), .Y95(Y95),
    .X96(X96), .Y96(Y96),
    .X97(X97), .Y97(Y97),
    .X98(X98), .Y98(Y98),
    .X99(X99), .Y99(Y99),
    .X100(X100), .Y100(Y100),
    .X101(X101), .Y101(Y101),
    .X102(X102), .Y102(Y102),
    .X103(X103), .Y103(Y103),
    .X104(X104), .Y104(Y104),
    .X105(X105), .Y105(Y105),
    .X106(X106), .Y106(Y106),
    .X107(X107), .Y107(Y107),
    .X108(X108), .Y108(Y108),
    .X109(X109), .Y109(Y109),
    .X110(X110), .Y110(Y110),
    .X111(X111), .Y111(Y111),
    .X112(X112), .Y112(Y112),
    .X113(X113), .Y113(Y113),
    .X114(X114), .Y114(Y114),
    .X115(X115), .Y115(Y115),
    .X116(X116), .Y116(Y116),
    .X117(X117), .Y117(Y117),
    .X118(X118), .Y118(Y118),
    .X119(X119), .Y119(Y119),
    .X120(X120), .Y120(Y120),
    .X121(X121), .Y121(Y121),
    .X122(X122), .Y122(Y122),
    .X123(X123), .Y123(Y123),
    .X124(X124), .Y124(Y124),
    .X125(X125), .Y125(Y125),
    .X126(X126), .Y126(Y126),
    .X127(X127), .Y127(Y127),
    .X128(X128), .Y128(Y128),
    .X129(X129), .Y129(Y129),
    .X130(X130), .Y130(Y130),
    .X131(X131), .Y131(Y131),
    .X132(X132), .Y132(Y132),
    .X133(X133), .Y133(Y133),
    .X134(X134), .Y134(Y134),
    .X135(X135), .Y135(Y135),
    .X136(X136), .Y136(Y136),
    .X137(X137), .Y137(Y137),
    .X138(X138), .Y138(Y138),
    .X139(X139), .Y139(Y139),
    .X140(X140), .Y140(Y140),
    .X141(X141), .Y141(Y141),
    .X142(X142), .Y142(Y142),
    .X143(X143), .Y143(Y143),
    .X144(X144), .Y144(Y144),
    .X145(X145), .Y145(Y145),
    .X146(X146), .Y146(Y146),
    .X147(X147), .Y147(Y147),
    .X148(X148), .Y148(Y148),
    .X149(X149), .Y149(Y149),
    .X150(X150), .Y150(Y150),
    .X151(X151), .Y151(Y151),
    .X152(X152), .Y152(Y152),
    .X153(X153), .Y153(Y153),
    .X154(X154), .Y154(Y154),
    .X155(X155), .Y155(Y155),
    .X156(X156), .Y156(Y156),
    .X157(X157), .Y157(Y157),
    .X158(X158), .Y158(Y158),
    .X159(X159), .Y159(Y159),
    .X160(X160), .Y160(Y160),
    .X161(X161), .Y161(Y161),
    .X162(X162), .Y162(Y162),
    .X163(X163), .Y163(Y163),
    .X164(X164), .Y164(Y164),
    .X165(X165), .Y165(Y165),
    .X166(X166), .Y166(Y166),
    .X167(X167), .Y167(Y167),
    .X168(X168), .Y168(Y168),
    .X169(X169), .Y169(Y169),
    .X170(X170), .Y170(Y170),
    .X171(X171), .Y171(Y171),
    .X172(X172), .Y172(Y172),
    .X173(X173), .Y173(Y173),
    .X174(X174), .Y174(Y174),
    .X175(X175), .Y175(Y175),
    .X176(X176), .Y176(Y176),
    .X177(X177), .Y177(Y177),
    .X178(X178), .Y178(Y178),
    .X179(X179), .Y179(Y179),
    .X180(X180), .Y180(Y180),
    .X181(X181), .Y181(Y181),
    .X182(X182), .Y182(Y182),
    .X183(X183), .Y183(Y183),
    .X184(X184), .Y184(Y184),
    .X185(X185), .Y185(Y185),
    .X186(X186), .Y186(Y186),
    .X187(X187), .Y187(Y187),
    .X188(X188), .Y188(Y188),
    .X189(X189), .Y189(Y189),
    .X190(X190), .Y190(Y190),
    .X191(X191), .Y191(Y191),
    .X192(X192), .Y192(Y192),
    .X193(X193), .Y193(Y193),
    .X194(X194), .Y194(Y194),
    .X195(X195), .Y195(Y195),
    .X196(X196), .Y196(Y196),
    .X197(X197), .Y197(Y197),
    .X198(X198), .Y198(Y198),
    .X199(X199), .Y199(Y199),
    .X200(X200), .Y200(Y200),
    .X201(X201), .Y201(Y201),
    .X202(X202), .Y202(Y202),
    .X203(X203), .Y203(Y203),
    .X204(X204), .Y204(Y204),
    .X205(X205), .Y205(Y205),
    .X206(X206), .Y206(Y206),
    .X207(X207), .Y207(Y207),
    .X208(X208), .Y208(Y208),
    .X209(X209), .Y209(Y209),
    .X210(X210), .Y210(Y210),
    .X211(X211), .Y211(Y211),
    .X212(X212), .Y212(Y212),
    .X213(X213), .Y213(Y213),
    .X214(X214), .Y214(Y214),
    .X215(X215), .Y215(Y215),
    .X216(X216), .Y216(Y216),
    .X217(X217), .Y217(Y217),
    .X218(X218), .Y218(Y218),
    .X219(X219), .Y219(Y219),
    .X220(X220), .Y220(Y220),
    .X221(X221), .Y221(Y221),
    .X222(X222), .Y222(Y222),
    .X223(X223), .Y223(Y223),
    .X224(X224), .Y224(Y224),
    .X225(X225), .Y225(Y225),
    .X226(X226), .Y226(Y226),
    .X227(X227), .Y227(Y227),
    .X228(X228), .Y228(Y228),
    .X229(X229), .Y229(Y229),
    .X230(X230), .Y230(Y230),
    .X231(X231), .Y231(Y231),
    .X232(X232), .Y232(Y232),
    .X233(X233), .Y233(Y233),
    .X234(X234), .Y234(Y234),
    .X235(X235), .Y235(Y235),
    .X236(X236), .Y236(Y236),
    .X237(X237), .Y237(Y237),
    .X238(X238), .Y238(Y238),
    .X239(X239), .Y239(Y239),
    .X240(X240), .Y240(Y240),
    .X241(X241), .Y241(Y241),
    .X242(X242), .Y242(Y242),
    .X243(X243), .Y243(Y243),
    .X244(X244), .Y244(Y244),
    .X245(X245), .Y245(Y245),
    .X246(X246), .Y246(Y246),
    .X247(X247), .Y247(Y247),
    .X248(X248), .Y248(Y248),
    .X249(X249), .Y249(Y249),
    .X250(X250), .Y250(Y250),
    .X251(X251), .Y251(Y251),
    .X252(X252), .Y252(Y252),
    .X253(X253), .Y253(Y253),
    .X254(X254), .Y254(Y254),
    .X255(X255), .Y255(Y255),
    .X256(X256), .Y256(Y256),
    .X257(X257), .Y257(Y257),
    .X258(X258), .Y258(Y258),
    .X259(X259), .Y259(Y259),
    .X260(X260), .Y260(Y260),
    .X261(X261), .Y261(Y261),
    .X262(X262), .Y262(Y262),
    .X263(X263), .Y263(Y263),
    .X264(X264), .Y264(Y264),
    .X265(X265), .Y265(Y265),
    .X266(X266), .Y266(Y266),
    .X267(X267), .Y267(Y267),
    .X268(X268), .Y268(Y268),
    .X269(X269), .Y269(Y269),
    .X270(X270), .Y270(Y270),
    .X271(X271), .Y271(Y271),
    .X272(X272), .Y272(Y272),
    .X273(X273), .Y273(Y273),
    .X274(X274), .Y274(Y274),
    .X275(X275), .Y275(Y275),
    .X276(X276), .Y276(Y276),
    .X277(X277), .Y277(Y277),
    .X278(X278), .Y278(Y278),
    .X279(X279), .Y279(Y279),
    .X280(X280), .Y280(Y280),
    .X281(X281), .Y281(Y281),
    .X282(X282), .Y282(Y282),
    .X283(X283), .Y283(Y283),
    .X284(X284), .Y284(Y284),
    .X285(X285), .Y285(Y285),
    .X286(X286), .Y286(Y286),
    .X287(X287), .Y287(Y287),
    .X288(X288), .Y288(Y288),
    .X289(X289), .Y289(Y289),
    .X290(X290), .Y290(Y290),
    .X291(X291), .Y291(Y291),
    .X292(X292), .Y292(Y292),
    .X293(X293), .Y293(Y293),
    .X294(X294), .Y294(Y294),
    .X295(X295), .Y295(Y295),
    .X296(X296), .Y296(Y296),
    .X297(X297), .Y297(Y297),
    .X298(X298), .Y298(Y298),
    .X299(X299), .Y299(Y299),
    .X300(X300), .Y300(Y300),
    .X301(X301), .Y301(Y301),
    .X302(X302), .Y302(Y302),
    .X303(X303), .Y303(Y303),
    .X304(X304), .Y304(Y304),
    .X305(X305), .Y305(Y305),
    .X306(X306), .Y306(Y306),
    .X307(X307), .Y307(Y307),
    .X308(X308), .Y308(Y308),
    .X309(X309), .Y309(Y309),
    .X310(X310), .Y310(Y310),
    .X311(X311), .Y311(Y311),
    .X312(X312), .Y312(Y312),
    .X313(X313), .Y313(Y313),
    .X314(X314), .Y314(Y314),
    .X315(X315), .Y315(Y315),
    .X316(X316), .Y316(Y316),
    .X317(X317), .Y317(Y317),
    .X318(X318), .Y318(Y318),
    .X319(X319), .Y319(Y319),
    .X320(X320), .Y320(Y320),
    .X321(X321), .Y321(Y321),
    .X322(X322), .Y322(Y322),
    .X323(X323), .Y323(Y323),
    .X324(X324), .Y324(Y324),
    .X325(X325), .Y325(Y325),
    .X326(X326), .Y326(Y326),
    .X327(X327), .Y327(Y327),
    .X328(X328), .Y328(Y328),
    .X329(X329), .Y329(Y329),
    .X330(X330), .Y330(Y330),
    .X331(X331), .Y331(Y331),
    .X332(X332), .Y332(Y332),
    .X333(X333), .Y333(Y333),
    .X334(X334), .Y334(Y334),
    .X335(X335), .Y335(Y335),
    .X336(X336), .Y336(Y336),
    .X337(X337), .Y337(Y337),
    .X338(X338), .Y338(Y338),
    .X339(X339), .Y339(Y339),
    .X340(X340), .Y340(Y340),
    .X341(X341), .Y341(Y341),
    .X342(X342), .Y342(Y342),
    .X343(X343), .Y343(Y343),
    .X344(X344), .Y344(Y344),
    .X345(X345), .Y345(Y345),
    .X346(X346), .Y346(Y346),
    .X347(X347), .Y347(Y347),
    .X348(X348), .Y348(Y348),
    .X349(X349), .Y349(Y349),
    .X350(X350), .Y350(Y350),
    .X351(X351), .Y351(Y351),
    .X352(X352), .Y352(Y352),
    .X353(X353), .Y353(Y353),
    .X354(X354), .Y354(Y354),
    .X355(X355), .Y355(Y355),
    .X356(X356), .Y356(Y356),
    .X357(X357), .Y357(Y357),
    .X358(X358), .Y358(Y358),
    .X359(X359), .Y359(Y359),
    .X360(X360), .Y360(Y360),
    .X361(X361), .Y361(Y361),
    .X362(X362), .Y362(Y362),
    .X363(X363), .Y363(Y363),
    .X364(X364), .Y364(Y364),
    .X365(X365), .Y365(Y365),
    .X366(X366), .Y366(Y366),
    .X367(X367), .Y367(Y367),
    .X368(X368), .Y368(Y368),
    .X369(X369), .Y369(Y369),
    .X370(X370), .Y370(Y370),
    .X371(X371), .Y371(Y371),
    .X372(X372), .Y372(Y372),
    .X373(X373), .Y373(Y373),
    .X374(X374), .Y374(Y374),
    .X375(X375), .Y375(Y375),
    .X376(X376), .Y376(Y376),
    .X377(X377), .Y377(Y377),
    .X378(X378), .Y378(Y378),
    .X379(X379), .Y379(Y379),
    .X380(X380), .Y380(Y380),
    .X381(X381), .Y381(Y381),
    .X382(X382), .Y382(Y382),
    .X383(X383), .Y383(Y383),
    .X384(X384), .Y384(Y384),
    .X385(X385), .Y385(Y385),
    .X386(X386), .Y386(Y386),
    .X387(X387), .Y387(Y387),
    .X388(X388), .Y388(Y388),
    .X389(X389), .Y389(Y389),
    .X390(X390), .Y390(Y390),
    .X391(X391), .Y391(Y391),
    .X392(X392), .Y392(Y392),
    .X393(X393), .Y393(Y393),
    .X394(X394), .Y394(Y394),
    .X395(X395), .Y395(Y395),
    .X396(X396), .Y396(Y396),
    .X397(X397), .Y397(Y397),
    .X398(X398), .Y398(Y398),
    .X399(X399), .Y399(Y399),
    .X400(X400), .Y400(Y400),
    .X401(X401), .Y401(Y401),
    .X402(X402), .Y402(Y402),
    .X403(X403), .Y403(Y403),
    .X404(X404), .Y404(Y404),
    .X405(X405), .Y405(Y405),
    .X406(X406), .Y406(Y406),
    .X407(X407), .Y407(Y407),
    .X408(X408), .Y408(Y408),
    .X409(X409), .Y409(Y409),
    .X410(X410), .Y410(Y410),
    .X411(X411), .Y411(Y411),
    .X412(X412), .Y412(Y412),
    .X413(X413), .Y413(Y413),
    .X414(X414), .Y414(Y414),
    .X415(X415), .Y415(Y415),
    .X416(X416), .Y416(Y416),
    .X417(X417), .Y417(Y417),
    .X418(X418), .Y418(Y418),
    .X419(X419), .Y419(Y419),
    .X420(X420), .Y420(Y420),
    .X421(X421), .Y421(Y421),
    .X422(X422), .Y422(Y422),
    .X423(X423), .Y423(Y423),
    .X424(X424), .Y424(Y424),
    .X425(X425), .Y425(Y425),
    .X426(X426), .Y426(Y426),
    .X427(X427), .Y427(Y427),
    .X428(X428), .Y428(Y428),
    .X429(X429), .Y429(Y429),
    .X430(X430), .Y430(Y430),
    .X431(X431), .Y431(Y431),
    .X432(X432), .Y432(Y432),
    .X433(X433), .Y433(Y433),
    .X434(X434), .Y434(Y434),
    .X435(X435), .Y435(Y435),
    .X436(X436), .Y436(Y436),
    .X437(X437), .Y437(Y437),
    .X438(X438), .Y438(Y438),
    .X439(X439), .Y439(Y439),
    .X440(X440), .Y440(Y440),
    .X441(X441), .Y441(Y441),
    .X442(X442), .Y442(Y442),
    .X443(X443), .Y443(Y443),
    .X444(X444), .Y444(Y444),
    .X445(X445), .Y445(Y445),
    .X446(X446), .Y446(Y446),
    .X447(X447), .Y447(Y447),
    .X448(X448), .Y448(Y448),
    .X449(X449), .Y449(Y449),
    .X450(X450), .Y450(Y450),
    .X451(X451), .Y451(Y451),
    .X452(X452), .Y452(Y452),
    .X453(X453), .Y453(Y453),
    .X454(X454), .Y454(Y454),
    .X455(X455), .Y455(Y455),
    .X456(X456), .Y456(Y456),
    .X457(X457), .Y457(Y457),
    .X458(X458), .Y458(Y458),
    .X459(X459), .Y459(Y459),
    .X460(X460), .Y460(Y460),
    .X461(X461), .Y461(Y461),
    .X462(X462), .Y462(Y462),
    .X463(X463), .Y463(Y463),
    .X464(X464), .Y464(Y464),
    .X465(X465), .Y465(Y465),
    .X466(X466), .Y466(Y466),
    .X467(X467), .Y467(Y467),
    .X468(X468), .Y468(Y468),
    .X469(X469), .Y469(Y469),
    .X470(X470), .Y470(Y470),
    .X471(X471), .Y471(Y471),
    .X472(X472), .Y472(Y472),
    .X473(X473), .Y473(Y473),
    .X474(X474), .Y474(Y474),
    .X475(X475), .Y475(Y475),
    .X476(X476), .Y476(Y476),
    .X477(X477), .Y477(Y477),
    .X478(X478), .Y478(Y478),
    .X479(X479), .Y479(Y479),
    .X480(X480), .Y480(Y480),
    .X481(X481), .Y481(Y481),
    .X482(X482), .Y482(Y482),
    .X483(X483), .Y483(Y483),
    .X484(X484), .Y484(Y484),
    .X485(X485), .Y485(Y485),
    .X486(X486), .Y486(Y486),
    .X487(X487), .Y487(Y487),
    .X488(X488), .Y488(Y488),
    .X489(X489), .Y489(Y489),
    .X490(X490), .Y490(Y490),
    .X491(X491), .Y491(Y491),
    .X492(X492), .Y492(Y492),
    .X493(X493), .Y493(Y493),
    .X494(X494), .Y494(Y494),
    .X495(X495), .Y495(Y495),
    .X496(X496), .Y496(Y496),
    .X497(X497), .Y497(Y497),
    .X498(X498), .Y498(Y498),
    .X499(X499), .Y499(Y499),
    .X500(X500), .Y500(Y500),
    .X501(X501), .Y501(Y501),
    .X502(X502), .Y502(Y502),
    .X503(X503), .Y503(Y503),
    .X504(X504), .Y504(Y504),
    .X505(X505), .Y505(Y505),
    .X506(X506), .Y506(Y506),
    .X507(X507), .Y507(Y507),
    .X508(X508), .Y508(Y508),
    .X509(X509), .Y509(Y509),
    .X510(X510), .Y510(Y510),
    .X511(X511), .Y511(Y511),
    .X512(X512), .Y512(Y512),
    .X513(X513), .Y513(Y513),
    .X514(X514), .Y514(Y514),
    .X515(X515), .Y515(Y515),
    .X516(X516), .Y516(Y516),
    .X517(X517), .Y517(Y517),
    .X518(X518), .Y518(Y518),
    .X519(X519), .Y519(Y519),
    .X520(X520), .Y520(Y520),
    .X521(X521), .Y521(Y521),
    .X522(X522), .Y522(Y522),
    .X523(X523), .Y523(Y523),
    .X524(X524), .Y524(Y524),
    .X525(X525), .Y525(Y525),
    .X526(X526), .Y526(Y526),
    .X527(X527), .Y527(Y527),
    .X528(X528), .Y528(Y528),
    .X529(X529), .Y529(Y529),
    .X530(X530), .Y530(Y530),
    .X531(X531), .Y531(Y531),
    .X532(X532), .Y532(Y532),
    .X533(X533), .Y533(Y533),
    .X534(X534), .Y534(Y534),
    .X535(X535), .Y535(Y535),
    .X536(X536), .Y536(Y536),
    .X537(X537), .Y537(Y537),
    .X538(X538), .Y538(Y538),
    .X539(X539), .Y539(Y539),
    .X540(X540), .Y540(Y540),
    .X541(X541), .Y541(Y541),
    .X542(X542), .Y542(Y542),
    .X543(X543), .Y543(Y543),
    .X544(X544), .Y544(Y544),
    .X545(X545), .Y545(Y545),
    .X546(X546), .Y546(Y546),
    .X547(X547), .Y547(Y547),
    .X548(X548), .Y548(Y548),
    .X549(X549), .Y549(Y549),
    .X550(X550), .Y550(Y550),
    .X551(X551), .Y551(Y551),
    .X552(X552), .Y552(Y552),
    .X553(X553), .Y553(Y553),
    .X554(X554), .Y554(Y554),
    .X555(X555), .Y555(Y555),
    .X556(X556), .Y556(Y556),
    .X557(X557), .Y557(Y557),
    .X558(X558), .Y558(Y558),
    .X559(X559), .Y559(Y559),
    .X560(X560), .Y560(Y560),
    .X561(X561), .Y561(Y561),
    .X562(X562), .Y562(Y562),
    .X563(X563), .Y563(Y563),
    .X564(X564), .Y564(Y564),
    .X565(X565), .Y565(Y565),
    .X566(X566), .Y566(Y566),
    .X567(X567), .Y567(Y567),
    .X568(X568), .Y568(Y568),
    .X569(X569), .Y569(Y569),
    .X570(X570), .Y570(Y570),
    .X571(X571), .Y571(Y571),
    .X572(X572), .Y572(Y572),
    .X573(X573), .Y573(Y573),
    .X574(X574), .Y574(Y574),
    .X575(X575), .Y575(Y575),
    .X576(X576), .Y576(Y576),
    .X577(X577), .Y577(Y577),
    .X578(X578), .Y578(Y578),
    .X579(X579), .Y579(Y579),
    .X580(X580), .Y580(Y580),
    .X581(X581), .Y581(Y581),
    .X582(X582), .Y582(Y582),
    .X583(X583), .Y583(Y583),
    .X584(X584), .Y584(Y584),
    .X585(X585), .Y585(Y585),
    .X586(X586), .Y586(Y586),
    .X587(X587), .Y587(Y587),
    .X588(X588), .Y588(Y588),
    .X589(X589), .Y589(Y589),
    .X590(X590), .Y590(Y590),
    .X591(X591), .Y591(Y591),
    .X592(X592), .Y592(Y592),
    .X593(X593), .Y593(Y593),
    .X594(X594), .Y594(Y594),
    .X595(X595), .Y595(Y595),
    .X596(X596), .Y596(Y596),
    .X597(X597), .Y597(Y597),
    .X598(X598), .Y598(Y598),
    .X599(X599), .Y599(Y599),
    .X600(X600), .Y600(Y600),
    .X601(X601), .Y601(Y601),
    .X602(X602), .Y602(Y602),
    .X603(X603), .Y603(Y603),
    .X604(X604), .Y604(Y604),
    .X605(X605), .Y605(Y605),
    .X606(X606), .Y606(Y606),
    .X607(X607), .Y607(Y607),
    .X608(X608), .Y608(Y608),
    .X609(X609), .Y609(Y609),
    .X610(X610), .Y610(Y610),
    .X611(X611), .Y611(Y611),
    .X612(X612), .Y612(Y612),
    .X613(X613), .Y613(Y613),
    .X614(X614), .Y614(Y614),
    .X615(X615), .Y615(Y615),
    .X616(X616), .Y616(Y616),
    .X617(X617), .Y617(Y617),
    .X618(X618), .Y618(Y618),
    .X619(X619), .Y619(Y619),
    .X620(X620), .Y620(Y620),
    .X621(X621), .Y621(Y621),
    .X622(X622), .Y622(Y622),
    .X623(X623), .Y623(Y623),
    .X624(X624), .Y624(Y624),
    .X625(X625), .Y625(Y625),
    .X626(X626), .Y626(Y626),
    .X627(X627), .Y627(Y627),
    .X628(X628), .Y628(Y628),
    .X629(X629), .Y629(Y629),
    .X630(X630), .Y630(Y630),
    .X631(X631), .Y631(Y631),
    .X632(X632), .Y632(Y632),
    .X633(X633), .Y633(Y633),
    .X634(X634), .Y634(Y634),
    .X635(X635), .Y635(Y635),
    .X636(X636), .Y636(Y636),
    .X637(X637), .Y637(Y637),
    .X638(X638), .Y638(Y638),
    .X639(X639), .Y639(Y639),
    .X640(X640), .Y640(Y640),
    .X641(X641), .Y641(Y641),
    .X642(X642), .Y642(Y642),
    .X643(X643), .Y643(Y643),
    .X644(X644), .Y644(Y644),
    .X645(X645), .Y645(Y645),
    .X646(X646), .Y646(Y646),
    .X647(X647), .Y647(Y647),
    .X648(X648), .Y648(Y648),
    .X649(X649), .Y649(Y649),
    .X650(X650), .Y650(Y650),
    .X651(X651), .Y651(Y651),
    .X652(X652), .Y652(Y652),
    .X653(X653), .Y653(Y653),
    .X654(X654), .Y654(Y654),
    .X655(X655), .Y655(Y655),
    .X656(X656), .Y656(Y656),
    .X657(X657), .Y657(Y657),
    .X658(X658), .Y658(Y658),
    .X659(X659), .Y659(Y659),
    .X660(X660), .Y660(Y660),
    .X661(X661), .Y661(Y661),
    .X662(X662), .Y662(Y662),
    .X663(X663), .Y663(Y663),
    .X664(X664), .Y664(Y664),
    .X665(X665), .Y665(Y665),
    .X666(X666), .Y666(Y666),
    .X667(X667), .Y667(Y667),
    .X668(X668), .Y668(Y668),
    .X669(X669), .Y669(Y669),
    .X670(X670), .Y670(Y670),
    .X671(X671), .Y671(Y671),
    .X672(X672), .Y672(Y672),
    .X673(X673), .Y673(Y673),
    .X674(X674), .Y674(Y674),
    .X675(X675), .Y675(Y675),
    .X676(X676), .Y676(Y676),
    .X677(X677), .Y677(Y677),
    .X678(X678), .Y678(Y678),
    .X679(X679), .Y679(Y679),
    .X680(X680), .Y680(Y680),
    .X681(X681), .Y681(Y681),
    .X682(X682), .Y682(Y682),
    .X683(X683), .Y683(Y683),
    .X684(X684), .Y684(Y684),
    .X685(X685), .Y685(Y685),
    .X686(X686), .Y686(Y686),
    .X687(X687), .Y687(Y687),
    .X688(X688), .Y688(Y688),
    .X689(X689), .Y689(Y689),
    .X690(X690), .Y690(Y690),
    .X691(X691), .Y691(Y691),
    .X692(X692), .Y692(Y692),
    .X693(X693), .Y693(Y693),
    .X694(X694), .Y694(Y694),
    .X695(X695), .Y695(Y695),
    .X696(X696), .Y696(Y696),
    .X697(X697), .Y697(Y697),
    .X698(X698), .Y698(Y698),
    .X699(X699), .Y699(Y699),
    .X700(X700), .Y700(Y700),
    .X701(X701), .Y701(Y701),
    .X702(X702), .Y702(Y702),
    .X703(X703), .Y703(Y703),
    .X704(X704), .Y704(Y704),
    .X705(X705), .Y705(Y705),
    .X706(X706), .Y706(Y706),
    .X707(X707), .Y707(Y707),
    .X708(X708), .Y708(Y708),
    .X709(X709), .Y709(Y709),
    .X710(X710), .Y710(Y710),
    .X711(X711), .Y711(Y711),
    .X712(X712), .Y712(Y712),
    .X713(X713), .Y713(Y713),
    .X714(X714), .Y714(Y714),
    .X715(X715), .Y715(Y715),
    .X716(X716), .Y716(Y716),
    .X717(X717), .Y717(Y717),
    .X718(X718), .Y718(Y718),
    .X719(X719), .Y719(Y719),
    .X720(X720), .Y720(Y720),
    .X721(X721), .Y721(Y721),
    .X722(X722), .Y722(Y722),
    .X723(X723), .Y723(Y723),
    .X724(X724), .Y724(Y724),
    .X725(X725), .Y725(Y725),
    .X726(X726), .Y726(Y726),
    .X727(X727), .Y727(Y727),
    .X728(X728), .Y728(Y728),
    .X729(X729), .Y729(Y729),
    .X730(X730), .Y730(Y730),
    .X731(X731), .Y731(Y731),
    .X732(X732), .Y732(Y732),
    .X733(X733), .Y733(Y733),
    .X734(X734), .Y734(Y734),
    .X735(X735), .Y735(Y735),
    .X736(X736), .Y736(Y736),
    .X737(X737), .Y737(Y737),
    .X738(X738), .Y738(Y738),
    .X739(X739), .Y739(Y739),
    .X740(X740), .Y740(Y740),
    .X741(X741), .Y741(Y741),
    .X742(X742), .Y742(Y742),
    .X743(X743), .Y743(Y743),
    .X744(X744), .Y744(Y744),
    .X745(X745), .Y745(Y745),
    .X746(X746), .Y746(Y746),
    .X747(X747), .Y747(Y747),
    .X748(X748), .Y748(Y748),
    .X749(X749), .Y749(Y749),
    .X750(X750), .Y750(Y750),
    .X751(X751), .Y751(Y751),
    .X752(X752), .Y752(Y752),
    .X753(X753), .Y753(Y753),
    .X754(X754), .Y754(Y754),
    .X755(X755), .Y755(Y755),
    .X756(X756), .Y756(Y756),
    .X757(X757), .Y757(Y757),
    .X758(X758), .Y758(Y758),
    .X759(X759), .Y759(Y759),
    .X760(X760), .Y760(Y760),
    .X761(X761), .Y761(Y761),
    .X762(X762), .Y762(Y762),
    .X763(X763), .Y763(Y763),
    .X764(X764), .Y764(Y764),
    .X765(X765), .Y765(Y765),
    .X766(X766), .Y766(Y766),
    .X767(X767), .Y767(Y767),
    .X768(X768), .Y768(Y768),
    .X769(X769), .Y769(Y769),
    .X770(X770), .Y770(Y770),
    .X771(X771), .Y771(Y771),
    .X772(X772), .Y772(Y772),
    .X773(X773), .Y773(Y773),
    .X774(X774), .Y774(Y774),
    .X775(X775), .Y775(Y775),
    .X776(X776), .Y776(Y776),
    .X777(X777), .Y777(Y777),
    .X778(X778), .Y778(Y778),
    .X779(X779), .Y779(Y779),
    .X780(X780), .Y780(Y780),
    .X781(X781), .Y781(Y781),
    .X782(X782), .Y782(Y782),
    .X783(X783), .Y783(Y783),
    .X784(X784), .Y784(Y784),
    .X785(X785), .Y785(Y785),
    .X786(X786), .Y786(Y786),
    .X787(X787), .Y787(Y787),
    .X788(X788), .Y788(Y788),
    .X789(X789), .Y789(Y789),
    .X790(X790), .Y790(Y790),
    .X791(X791), .Y791(Y791),
    .X792(X792), .Y792(Y792),
    .X793(X793), .Y793(Y793),
    .X794(X794), .Y794(Y794),
    .X795(X795), .Y795(Y795),
    .X796(X796), .Y796(Y796),
    .X797(X797), .Y797(Y797),
    .X798(X798), .Y798(Y798),
    .X799(X799), .Y799(Y799),
    .X800(X800), .Y800(Y800),
    .X801(X801), .Y801(Y801),
    .X802(X802), .Y802(Y802),
    .X803(X803), .Y803(Y803),
    .X804(X804), .Y804(Y804),
    .X805(X805), .Y805(Y805),
    .X806(X806), .Y806(Y806),
    .X807(X807), .Y807(Y807),
    .X808(X808), .Y808(Y808),
    .X809(X809), .Y809(Y809),
    .X810(X810), .Y810(Y810),
    .X811(X811), .Y811(Y811),
    .X812(X812), .Y812(Y812),
    .X813(X813), .Y813(Y813),
    .X814(X814), .Y814(Y814),
    .X815(X815), .Y815(Y815),
    .X816(X816), .Y816(Y816),
    .X817(X817), .Y817(Y817),
    .X818(X818), .Y818(Y818),
    .X819(X819), .Y819(Y819),
    .X820(X820), .Y820(Y820),
    .X821(X821), .Y821(Y821),
    .X822(X822), .Y822(Y822),
    .X823(X823), .Y823(Y823),
    .X824(X824), .Y824(Y824),
    .X825(X825), .Y825(Y825),
    .X826(X826), .Y826(Y826),
    .X827(X827), .Y827(Y827),
    .X828(X828), .Y828(Y828),
    .X829(X829), .Y829(Y829),
    .X830(X830), .Y830(Y830),
    .X831(X831), .Y831(Y831),
    .X832(X832), .Y832(Y832),
    .X833(X833), .Y833(Y833),
    .X834(X834), .Y834(Y834),
    .X835(X835), .Y835(Y835),
    .X836(X836), .Y836(Y836),
    .X837(X837), .Y837(Y837),
    .X838(X838), .Y838(Y838),
    .X839(X839), .Y839(Y839),
    .X840(X840), .Y840(Y840),
    .X841(X841), .Y841(Y841),
    .X842(X842), .Y842(Y842),
    .X843(X843), .Y843(Y843),
    .X844(X844), .Y844(Y844),
    .X845(X845), .Y845(Y845),
    .X846(X846), .Y846(Y846),
    .X847(X847), .Y847(Y847),
    .X848(X848), .Y848(Y848),
    .X849(X849), .Y849(Y849),
    .X850(X850), .Y850(Y850),
    .X851(X851), .Y851(Y851),
    .X852(X852), .Y852(Y852),
    .X853(X853), .Y853(Y853),
    .X854(X854), .Y854(Y854),
    .X855(X855), .Y855(Y855),
    .X856(X856), .Y856(Y856),
    .X857(X857), .Y857(Y857),
    .X858(X858), .Y858(Y858),
    .X859(X859), .Y859(Y859),
    .X860(X860), .Y860(Y860),
    .X861(X861), .Y861(Y861),
    .X862(X862), .Y862(Y862),
    .X863(X863), .Y863(Y863),
    .X864(X864), .Y864(Y864),
    .X865(X865), .Y865(Y865),
    .X866(X866), .Y866(Y866),
    .X867(X867), .Y867(Y867),
    .X868(X868), .Y868(Y868),
    .X869(X869), .Y869(Y869),
    .X870(X870), .Y870(Y870),
    .X871(X871), .Y871(Y871),
    .X872(X872), .Y872(Y872),
    .X873(X873), .Y873(Y873),
    .X874(X874), .Y874(Y874),
    .X875(X875), .Y875(Y875),
    .X876(X876), .Y876(Y876),
    .X877(X877), .Y877(Y877),
    .X878(X878), .Y878(Y878),
    .X879(X879), .Y879(Y879),
    .X880(X880), .Y880(Y880),
    .X881(X881), .Y881(Y881),
    .X882(X882), .Y882(Y882),
    .X883(X883), .Y883(Y883),
    .X884(X884), .Y884(Y884),
    .X885(X885), .Y885(Y885),
    .X886(X886), .Y886(Y886),
    .X887(X887), .Y887(Y887),
    .X888(X888), .Y888(Y888),
    .X889(X889), .Y889(Y889),
    .X890(X890), .Y890(Y890),
    .X891(X891), .Y891(Y891),
    .X892(X892), .Y892(Y892),
    .X893(X893), .Y893(Y893),
    .X894(X894), .Y894(Y894),
    .X895(X895), .Y895(Y895),
    .X896(X896), .Y896(Y896),
    .X897(X897), .Y897(Y897),
    .X898(X898), .Y898(Y898),
    .X899(X899), .Y899(Y899),
    .X900(X900), .Y900(Y900),
    .X901(X901), .Y901(Y901),
    .X902(X902), .Y902(Y902),
    .X903(X903), .Y903(Y903),
    .X904(X904), .Y904(Y904),
    .X905(X905), .Y905(Y905),
    .X906(X906), .Y906(Y906),
    .X907(X907), .Y907(Y907),
    .X908(X908), .Y908(Y908),
    .X909(X909), .Y909(Y909),
    .X910(X910), .Y910(Y910),
    .X911(X911), .Y911(Y911),
    .X912(X912), .Y912(Y912),
    .X913(X913), .Y913(Y913),
    .X914(X914), .Y914(Y914),
    .X915(X915), .Y915(Y915),
    .X916(X916), .Y916(Y916),
    .X917(X917), .Y917(Y917),
    .X918(X918), .Y918(Y918),
    .X919(X919), .Y919(Y919),
    .X920(X920), .Y920(Y920),
    .X921(X921), .Y921(Y921),
    .X922(X922), .Y922(Y922),
    .X923(X923), .Y923(Y923),
    .X924(X924), .Y924(Y924),
    .X925(X925), .Y925(Y925),
    .X926(X926), .Y926(Y926),
    .X927(X927), .Y927(Y927),
    .X928(X928), .Y928(Y928),
    .X929(X929), .Y929(Y929),
    .X930(X930), .Y930(Y930),
    .X931(X931), .Y931(Y931),
    .X932(X932), .Y932(Y932),
    .X933(X933), .Y933(Y933),
    .X934(X934), .Y934(Y934),
    .X935(X935), .Y935(Y935),
    .X936(X936), .Y936(Y936),
    .X937(X937), .Y937(Y937),
    .X938(X938), .Y938(Y938),
    .X939(X939), .Y939(Y939),
    .X940(X940), .Y940(Y940),
    .X941(X941), .Y941(Y941),
    .X942(X942), .Y942(Y942),
    .X943(X943), .Y943(Y943),
    .X944(X944), .Y944(Y944),
    .X945(X945), .Y945(Y945),
    .X946(X946), .Y946(Y946),
    .X947(X947), .Y947(Y947),
    .X948(X948), .Y948(Y948),
    .X949(X949), .Y949(Y949),
    .X950(X950), .Y950(Y950),
    .X951(X951), .Y951(Y951),
    .X952(X952), .Y952(Y952),
    .X953(X953), .Y953(Y953),
    .X954(X954), .Y954(Y954),
    .X955(X955), .Y955(Y955),
    .X956(X956), .Y956(Y956),
    .X957(X957), .Y957(Y957),
    .X958(X958), .Y958(Y958),
    .X959(X959), .Y959(Y959),
    .X960(X960), .Y960(Y960),
    .X961(X961), .Y961(Y961),
    .X962(X962), .Y962(Y962),
    .X963(X963), .Y963(Y963),
    .X964(X964), .Y964(Y964),
    .X965(X965), .Y965(Y965),
    .X966(X966), .Y966(Y966),
    .X967(X967), .Y967(Y967),
    .X968(X968), .Y968(Y968),
    .X969(X969), .Y969(Y969),
    .X970(X970), .Y970(Y970),
    .X971(X971), .Y971(Y971),
    .X972(X972), .Y972(Y972),
    .X973(X973), .Y973(Y973),
    .X974(X974), .Y974(Y974),
    .X975(X975), .Y975(Y975),
    .X976(X976), .Y976(Y976),
    .X977(X977), .Y977(Y977),
    .X978(X978), .Y978(Y978),
    .X979(X979), .Y979(Y979),
    .X980(X980), .Y980(Y980),
    .X981(X981), .Y981(Y981),
    .X982(X982), .Y982(Y982),
    .X983(X983), .Y983(Y983),
    .X984(X984), .Y984(Y984),
    .X985(X985), .Y985(Y985),
    .X986(X986), .Y986(Y986),
    .X987(X987), .Y987(Y987),
    .X988(X988), .Y988(Y988),
    .X989(X989), .Y989(Y989),
    .X990(X990), .Y990(Y990),
    .X991(X991), .Y991(Y991),
    .X992(X992), .Y992(Y992),
    .X993(X993), .Y993(Y993),
    .X994(X994), .Y994(Y994),
    .X995(X995), .Y995(Y995),
    .X996(X996), .Y996(Y996),
    .X997(X997), .Y997(Y997),
    .X998(X998), .Y998(Y998),
    .X999(X999), .Y999(Y999),
    .X1000(X1000), .Y1000(Y1000),
    .X1001(X1001), .Y1001(Y1001),
    .X1002(X1002), .Y1002(Y1002),
    .X1003(X1003), .Y1003(Y1003),
    .X1004(X1004), .Y1004(Y1004),
    .X1005(X1005), .Y1005(Y1005),
    .X1006(X1006), .Y1006(Y1006),
    .X1007(X1007), .Y1007(Y1007),
    .X1008(X1008), .Y1008(Y1008),
    .X1009(X1009), .Y1009(Y1009),
    .X1010(X1010), .Y1010(Y1010),
    .X1011(X1011), .Y1011(Y1011),
    .X1012(X1012), .Y1012(Y1012),
    .X1013(X1013), .Y1013(Y1013),
    .X1014(X1014), .Y1014(Y1014),
    .X1015(X1015), .Y1015(Y1015),
    .X1016(X1016), .Y1016(Y1016),
    .X1017(X1017), .Y1017(Y1017),
    .X1018(X1018), .Y1018(Y1018),
    .X1019(X1019), .Y1019(Y1019),
    .X1020(X1020), .Y1020(Y1020),
    .X1021(X1021), .Y1021(Y1021),
    .X1022(X1022), .Y1022(Y1022),
    .X1023(X1023), .Y1023(Y1023));

   // You can use this counter to verify that the gap and latency are as expected.
   always @(posedge clk) begin
      if (clrCnt) counter <= 0;
      else counter <= counter+1;
   end


   initial begin
      @(posedge clk);
      @(posedge clk);

      // On the next cycle, begin loading input vector.
      next <= 1;
      clrCnt <= 1;
      @(posedge clk);
      clrCnt <= 0;
      next <= 0;

      // The 512 complex data points enter the system over 1 cycles
      for (j=0; j < 0; j = j+1) begin
          // Input: 512 complex words per cycle
         for (k=0; k < 1024; k = k+1) begin
            in[k] <= j*1024 + k;
         end
         @(posedge clk);
      end
      j = 0;
      for (k=0; k < 1024; k = k+1) begin
         in[k] <= j*1024 + k;
      end


      @(posedge clk);
      // Wait until the next data vector can be entered
      while (counter < 86)
        @(posedge clk);

      // On the next cycle, we will start the next data vector
      next <= 1;
      clrCnt <= 1;
      @(posedge clk);
      clrCnt <= 0;
      next <= 0;

      // Start entering next input vector
      for (j=0; j < 0; j = j+1) begin
         // Input 1024 words per cycle
         for (k=0; k < 1024; k = k+1) begin
            in[k] <= 1024 + j*1024 + k;
          end
          @(posedge clk);
       end
       j = 0;
       for (k=0; k < 1024; k = k+1) begin
          in[k] <= 1024 + j*1024 + k;
       end
   end


   initial begin
      // set initial values
      in[0] <= 0;
      in[1] <= 0;
      in[2] <= 0;
      in[3] <= 0;
      in[4] <= 0;
      in[5] <= 0;
      in[6] <= 0;
      in[7] <= 0;
      in[8] <= 0;
      in[9] <= 0;
      in[10] <= 0;
      in[11] <= 0;
      in[12] <= 0;
      in[13] <= 0;
      in[14] <= 0;
      in[15] <= 0;
      in[16] <= 0;
      in[17] <= 0;
      in[18] <= 0;
      in[19] <= 0;
      in[20] <= 0;
      in[21] <= 0;
      in[22] <= 0;
      in[23] <= 0;
      in[24] <= 0;
      in[25] <= 0;
      in[26] <= 0;
      in[27] <= 0;
      in[28] <= 0;
      in[29] <= 0;
      in[30] <= 0;
      in[31] <= 0;
      in[32] <= 0;
      in[33] <= 0;
      in[34] <= 0;
      in[35] <= 0;
      in[36] <= 0;
      in[37] <= 0;
      in[38] <= 0;
      in[39] <= 0;
      in[40] <= 0;
      in[41] <= 0;
      in[42] <= 0;
      in[43] <= 0;
      in[44] <= 0;
      in[45] <= 0;
      in[46] <= 0;
      in[47] <= 0;
      in[48] <= 0;
      in[49] <= 0;
      in[50] <= 0;
      in[51] <= 0;
      in[52] <= 0;
      in[53] <= 0;
      in[54] <= 0;
      in[55] <= 0;
      in[56] <= 0;
      in[57] <= 0;
      in[58] <= 0;
      in[59] <= 0;
      in[60] <= 0;
      in[61] <= 0;
      in[62] <= 0;
      in[63] <= 0;
      in[64] <= 0;
      in[65] <= 0;
      in[66] <= 0;
      in[67] <= 0;
      in[68] <= 0;
      in[69] <= 0;
      in[70] <= 0;
      in[71] <= 0;
      in[72] <= 0;
      in[73] <= 0;
      in[74] <= 0;
      in[75] <= 0;
      in[76] <= 0;
      in[77] <= 0;
      in[78] <= 0;
      in[79] <= 0;
      in[80] <= 0;
      in[81] <= 0;
      in[82] <= 0;
      in[83] <= 0;
      in[84] <= 0;
      in[85] <= 0;
      in[86] <= 0;
      in[87] <= 0;
      in[88] <= 0;
      in[89] <= 0;
      in[90] <= 0;
      in[91] <= 0;
      in[92] <= 0;
      in[93] <= 0;
      in[94] <= 0;
      in[95] <= 0;
      in[96] <= 0;
      in[97] <= 0;
      in[98] <= 0;
      in[99] <= 0;
      in[100] <= 0;
      in[101] <= 0;
      in[102] <= 0;
      in[103] <= 0;
      in[104] <= 0;
      in[105] <= 0;
      in[106] <= 0;
      in[107] <= 0;
      in[108] <= 0;
      in[109] <= 0;
      in[110] <= 0;
      in[111] <= 0;
      in[112] <= 0;
      in[113] <= 0;
      in[114] <= 0;
      in[115] <= 0;
      in[116] <= 0;
      in[117] <= 0;
      in[118] <= 0;
      in[119] <= 0;
      in[120] <= 0;
      in[121] <= 0;
      in[122] <= 0;
      in[123] <= 0;
      in[124] <= 0;
      in[125] <= 0;
      in[126] <= 0;
      in[127] <= 0;
      in[128] <= 0;
      in[129] <= 0;
      in[130] <= 0;
      in[131] <= 0;
      in[132] <= 0;
      in[133] <= 0;
      in[134] <= 0;
      in[135] <= 0;
      in[136] <= 0;
      in[137] <= 0;
      in[138] <= 0;
      in[139] <= 0;
      in[140] <= 0;
      in[141] <= 0;
      in[142] <= 0;
      in[143] <= 0;
      in[144] <= 0;
      in[145] <= 0;
      in[146] <= 0;
      in[147] <= 0;
      in[148] <= 0;
      in[149] <= 0;
      in[150] <= 0;
      in[151] <= 0;
      in[152] <= 0;
      in[153] <= 0;
      in[154] <= 0;
      in[155] <= 0;
      in[156] <= 0;
      in[157] <= 0;
      in[158] <= 0;
      in[159] <= 0;
      in[160] <= 0;
      in[161] <= 0;
      in[162] <= 0;
      in[163] <= 0;
      in[164] <= 0;
      in[165] <= 0;
      in[166] <= 0;
      in[167] <= 0;
      in[168] <= 0;
      in[169] <= 0;
      in[170] <= 0;
      in[171] <= 0;
      in[172] <= 0;
      in[173] <= 0;
      in[174] <= 0;
      in[175] <= 0;
      in[176] <= 0;
      in[177] <= 0;
      in[178] <= 0;
      in[179] <= 0;
      in[180] <= 0;
      in[181] <= 0;
      in[182] <= 0;
      in[183] <= 0;
      in[184] <= 0;
      in[185] <= 0;
      in[186] <= 0;
      in[187] <= 0;
      in[188] <= 0;
      in[189] <= 0;
      in[190] <= 0;
      in[191] <= 0;
      in[192] <= 0;
      in[193] <= 0;
      in[194] <= 0;
      in[195] <= 0;
      in[196] <= 0;
      in[197] <= 0;
      in[198] <= 0;
      in[199] <= 0;
      in[200] <= 0;
      in[201] <= 0;
      in[202] <= 0;
      in[203] <= 0;
      in[204] <= 0;
      in[205] <= 0;
      in[206] <= 0;
      in[207] <= 0;
      in[208] <= 0;
      in[209] <= 0;
      in[210] <= 0;
      in[211] <= 0;
      in[212] <= 0;
      in[213] <= 0;
      in[214] <= 0;
      in[215] <= 0;
      in[216] <= 0;
      in[217] <= 0;
      in[218] <= 0;
      in[219] <= 0;
      in[220] <= 0;
      in[221] <= 0;
      in[222] <= 0;
      in[223] <= 0;
      in[224] <= 0;
      in[225] <= 0;
      in[226] <= 0;
      in[227] <= 0;
      in[228] <= 0;
      in[229] <= 0;
      in[230] <= 0;
      in[231] <= 0;
      in[232] <= 0;
      in[233] <= 0;
      in[234] <= 0;
      in[235] <= 0;
      in[236] <= 0;
      in[237] <= 0;
      in[238] <= 0;
      in[239] <= 0;
      in[240] <= 0;
      in[241] <= 0;
      in[242] <= 0;
      in[243] <= 0;
      in[244] <= 0;
      in[245] <= 0;
      in[246] <= 0;
      in[247] <= 0;
      in[248] <= 0;
      in[249] <= 0;
      in[250] <= 0;
      in[251] <= 0;
      in[252] <= 0;
      in[253] <= 0;
      in[254] <= 0;
      in[255] <= 0;
      in[256] <= 0;
      in[257] <= 0;
      in[258] <= 0;
      in[259] <= 0;
      in[260] <= 0;
      in[261] <= 0;
      in[262] <= 0;
      in[263] <= 0;
      in[264] <= 0;
      in[265] <= 0;
      in[266] <= 0;
      in[267] <= 0;
      in[268] <= 0;
      in[269] <= 0;
      in[270] <= 0;
      in[271] <= 0;
      in[272] <= 0;
      in[273] <= 0;
      in[274] <= 0;
      in[275] <= 0;
      in[276] <= 0;
      in[277] <= 0;
      in[278] <= 0;
      in[279] <= 0;
      in[280] <= 0;
      in[281] <= 0;
      in[282] <= 0;
      in[283] <= 0;
      in[284] <= 0;
      in[285] <= 0;
      in[286] <= 0;
      in[287] <= 0;
      in[288] <= 0;
      in[289] <= 0;
      in[290] <= 0;
      in[291] <= 0;
      in[292] <= 0;
      in[293] <= 0;
      in[294] <= 0;
      in[295] <= 0;
      in[296] <= 0;
      in[297] <= 0;
      in[298] <= 0;
      in[299] <= 0;
      in[300] <= 0;
      in[301] <= 0;
      in[302] <= 0;
      in[303] <= 0;
      in[304] <= 0;
      in[305] <= 0;
      in[306] <= 0;
      in[307] <= 0;
      in[308] <= 0;
      in[309] <= 0;
      in[310] <= 0;
      in[311] <= 0;
      in[312] <= 0;
      in[313] <= 0;
      in[314] <= 0;
      in[315] <= 0;
      in[316] <= 0;
      in[317] <= 0;
      in[318] <= 0;
      in[319] <= 0;
      in[320] <= 0;
      in[321] <= 0;
      in[322] <= 0;
      in[323] <= 0;
      in[324] <= 0;
      in[325] <= 0;
      in[326] <= 0;
      in[327] <= 0;
      in[328] <= 0;
      in[329] <= 0;
      in[330] <= 0;
      in[331] <= 0;
      in[332] <= 0;
      in[333] <= 0;
      in[334] <= 0;
      in[335] <= 0;
      in[336] <= 0;
      in[337] <= 0;
      in[338] <= 0;
      in[339] <= 0;
      in[340] <= 0;
      in[341] <= 0;
      in[342] <= 0;
      in[343] <= 0;
      in[344] <= 0;
      in[345] <= 0;
      in[346] <= 0;
      in[347] <= 0;
      in[348] <= 0;
      in[349] <= 0;
      in[350] <= 0;
      in[351] <= 0;
      in[352] <= 0;
      in[353] <= 0;
      in[354] <= 0;
      in[355] <= 0;
      in[356] <= 0;
      in[357] <= 0;
      in[358] <= 0;
      in[359] <= 0;
      in[360] <= 0;
      in[361] <= 0;
      in[362] <= 0;
      in[363] <= 0;
      in[364] <= 0;
      in[365] <= 0;
      in[366] <= 0;
      in[367] <= 0;
      in[368] <= 0;
      in[369] <= 0;
      in[370] <= 0;
      in[371] <= 0;
      in[372] <= 0;
      in[373] <= 0;
      in[374] <= 0;
      in[375] <= 0;
      in[376] <= 0;
      in[377] <= 0;
      in[378] <= 0;
      in[379] <= 0;
      in[380] <= 0;
      in[381] <= 0;
      in[382] <= 0;
      in[383] <= 0;
      in[384] <= 0;
      in[385] <= 0;
      in[386] <= 0;
      in[387] <= 0;
      in[388] <= 0;
      in[389] <= 0;
      in[390] <= 0;
      in[391] <= 0;
      in[392] <= 0;
      in[393] <= 0;
      in[394] <= 0;
      in[395] <= 0;
      in[396] <= 0;
      in[397] <= 0;
      in[398] <= 0;
      in[399] <= 0;
      in[400] <= 0;
      in[401] <= 0;
      in[402] <= 0;
      in[403] <= 0;
      in[404] <= 0;
      in[405] <= 0;
      in[406] <= 0;
      in[407] <= 0;
      in[408] <= 0;
      in[409] <= 0;
      in[410] <= 0;
      in[411] <= 0;
      in[412] <= 0;
      in[413] <= 0;
      in[414] <= 0;
      in[415] <= 0;
      in[416] <= 0;
      in[417] <= 0;
      in[418] <= 0;
      in[419] <= 0;
      in[420] <= 0;
      in[421] <= 0;
      in[422] <= 0;
      in[423] <= 0;
      in[424] <= 0;
      in[425] <= 0;
      in[426] <= 0;
      in[427] <= 0;
      in[428] <= 0;
      in[429] <= 0;
      in[430] <= 0;
      in[431] <= 0;
      in[432] <= 0;
      in[433] <= 0;
      in[434] <= 0;
      in[435] <= 0;
      in[436] <= 0;
      in[437] <= 0;
      in[438] <= 0;
      in[439] <= 0;
      in[440] <= 0;
      in[441] <= 0;
      in[442] <= 0;
      in[443] <= 0;
      in[444] <= 0;
      in[445] <= 0;
      in[446] <= 0;
      in[447] <= 0;
      in[448] <= 0;
      in[449] <= 0;
      in[450] <= 0;
      in[451] <= 0;
      in[452] <= 0;
      in[453] <= 0;
      in[454] <= 0;
      in[455] <= 0;
      in[456] <= 0;
      in[457] <= 0;
      in[458] <= 0;
      in[459] <= 0;
      in[460] <= 0;
      in[461] <= 0;
      in[462] <= 0;
      in[463] <= 0;
      in[464] <= 0;
      in[465] <= 0;
      in[466] <= 0;
      in[467] <= 0;
      in[468] <= 0;
      in[469] <= 0;
      in[470] <= 0;
      in[471] <= 0;
      in[472] <= 0;
      in[473] <= 0;
      in[474] <= 0;
      in[475] <= 0;
      in[476] <= 0;
      in[477] <= 0;
      in[478] <= 0;
      in[479] <= 0;
      in[480] <= 0;
      in[481] <= 0;
      in[482] <= 0;
      in[483] <= 0;
      in[484] <= 0;
      in[485] <= 0;
      in[486] <= 0;
      in[487] <= 0;
      in[488] <= 0;
      in[489] <= 0;
      in[490] <= 0;
      in[491] <= 0;
      in[492] <= 0;
      in[493] <= 0;
      in[494] <= 0;
      in[495] <= 0;
      in[496] <= 0;
      in[497] <= 0;
      in[498] <= 0;
      in[499] <= 0;
      in[500] <= 0;
      in[501] <= 0;
      in[502] <= 0;
      in[503] <= 0;
      in[504] <= 0;
      in[505] <= 0;
      in[506] <= 0;
      in[507] <= 0;
      in[508] <= 0;
      in[509] <= 0;
      in[510] <= 0;
      in[511] <= 0;
      in[512] <= 0;
      in[513] <= 0;
      in[514] <= 0;
      in[515] <= 0;
      in[516] <= 0;
      in[517] <= 0;
      in[518] <= 0;
      in[519] <= 0;
      in[520] <= 0;
      in[521] <= 0;
      in[522] <= 0;
      in[523] <= 0;
      in[524] <= 0;
      in[525] <= 0;
      in[526] <= 0;
      in[527] <= 0;
      in[528] <= 0;
      in[529] <= 0;
      in[530] <= 0;
      in[531] <= 0;
      in[532] <= 0;
      in[533] <= 0;
      in[534] <= 0;
      in[535] <= 0;
      in[536] <= 0;
      in[537] <= 0;
      in[538] <= 0;
      in[539] <= 0;
      in[540] <= 0;
      in[541] <= 0;
      in[542] <= 0;
      in[543] <= 0;
      in[544] <= 0;
      in[545] <= 0;
      in[546] <= 0;
      in[547] <= 0;
      in[548] <= 0;
      in[549] <= 0;
      in[550] <= 0;
      in[551] <= 0;
      in[552] <= 0;
      in[553] <= 0;
      in[554] <= 0;
      in[555] <= 0;
      in[556] <= 0;
      in[557] <= 0;
      in[558] <= 0;
      in[559] <= 0;
      in[560] <= 0;
      in[561] <= 0;
      in[562] <= 0;
      in[563] <= 0;
      in[564] <= 0;
      in[565] <= 0;
      in[566] <= 0;
      in[567] <= 0;
      in[568] <= 0;
      in[569] <= 0;
      in[570] <= 0;
      in[571] <= 0;
      in[572] <= 0;
      in[573] <= 0;
      in[574] <= 0;
      in[575] <= 0;
      in[576] <= 0;
      in[577] <= 0;
      in[578] <= 0;
      in[579] <= 0;
      in[580] <= 0;
      in[581] <= 0;
      in[582] <= 0;
      in[583] <= 0;
      in[584] <= 0;
      in[585] <= 0;
      in[586] <= 0;
      in[587] <= 0;
      in[588] <= 0;
      in[589] <= 0;
      in[590] <= 0;
      in[591] <= 0;
      in[592] <= 0;
      in[593] <= 0;
      in[594] <= 0;
      in[595] <= 0;
      in[596] <= 0;
      in[597] <= 0;
      in[598] <= 0;
      in[599] <= 0;
      in[600] <= 0;
      in[601] <= 0;
      in[602] <= 0;
      in[603] <= 0;
      in[604] <= 0;
      in[605] <= 0;
      in[606] <= 0;
      in[607] <= 0;
      in[608] <= 0;
      in[609] <= 0;
      in[610] <= 0;
      in[611] <= 0;
      in[612] <= 0;
      in[613] <= 0;
      in[614] <= 0;
      in[615] <= 0;
      in[616] <= 0;
      in[617] <= 0;
      in[618] <= 0;
      in[619] <= 0;
      in[620] <= 0;
      in[621] <= 0;
      in[622] <= 0;
      in[623] <= 0;
      in[624] <= 0;
      in[625] <= 0;
      in[626] <= 0;
      in[627] <= 0;
      in[628] <= 0;
      in[629] <= 0;
      in[630] <= 0;
      in[631] <= 0;
      in[632] <= 0;
      in[633] <= 0;
      in[634] <= 0;
      in[635] <= 0;
      in[636] <= 0;
      in[637] <= 0;
      in[638] <= 0;
      in[639] <= 0;
      in[640] <= 0;
      in[641] <= 0;
      in[642] <= 0;
      in[643] <= 0;
      in[644] <= 0;
      in[645] <= 0;
      in[646] <= 0;
      in[647] <= 0;
      in[648] <= 0;
      in[649] <= 0;
      in[650] <= 0;
      in[651] <= 0;
      in[652] <= 0;
      in[653] <= 0;
      in[654] <= 0;
      in[655] <= 0;
      in[656] <= 0;
      in[657] <= 0;
      in[658] <= 0;
      in[659] <= 0;
      in[660] <= 0;
      in[661] <= 0;
      in[662] <= 0;
      in[663] <= 0;
      in[664] <= 0;
      in[665] <= 0;
      in[666] <= 0;
      in[667] <= 0;
      in[668] <= 0;
      in[669] <= 0;
      in[670] <= 0;
      in[671] <= 0;
      in[672] <= 0;
      in[673] <= 0;
      in[674] <= 0;
      in[675] <= 0;
      in[676] <= 0;
      in[677] <= 0;
      in[678] <= 0;
      in[679] <= 0;
      in[680] <= 0;
      in[681] <= 0;
      in[682] <= 0;
      in[683] <= 0;
      in[684] <= 0;
      in[685] <= 0;
      in[686] <= 0;
      in[687] <= 0;
      in[688] <= 0;
      in[689] <= 0;
      in[690] <= 0;
      in[691] <= 0;
      in[692] <= 0;
      in[693] <= 0;
      in[694] <= 0;
      in[695] <= 0;
      in[696] <= 0;
      in[697] <= 0;
      in[698] <= 0;
      in[699] <= 0;
      in[700] <= 0;
      in[701] <= 0;
      in[702] <= 0;
      in[703] <= 0;
      in[704] <= 0;
      in[705] <= 0;
      in[706] <= 0;
      in[707] <= 0;
      in[708] <= 0;
      in[709] <= 0;
      in[710] <= 0;
      in[711] <= 0;
      in[712] <= 0;
      in[713] <= 0;
      in[714] <= 0;
      in[715] <= 0;
      in[716] <= 0;
      in[717] <= 0;
      in[718] <= 0;
      in[719] <= 0;
      in[720] <= 0;
      in[721] <= 0;
      in[722] <= 0;
      in[723] <= 0;
      in[724] <= 0;
      in[725] <= 0;
      in[726] <= 0;
      in[727] <= 0;
      in[728] <= 0;
      in[729] <= 0;
      in[730] <= 0;
      in[731] <= 0;
      in[732] <= 0;
      in[733] <= 0;
      in[734] <= 0;
      in[735] <= 0;
      in[736] <= 0;
      in[737] <= 0;
      in[738] <= 0;
      in[739] <= 0;
      in[740] <= 0;
      in[741] <= 0;
      in[742] <= 0;
      in[743] <= 0;
      in[744] <= 0;
      in[745] <= 0;
      in[746] <= 0;
      in[747] <= 0;
      in[748] <= 0;
      in[749] <= 0;
      in[750] <= 0;
      in[751] <= 0;
      in[752] <= 0;
      in[753] <= 0;
      in[754] <= 0;
      in[755] <= 0;
      in[756] <= 0;
      in[757] <= 0;
      in[758] <= 0;
      in[759] <= 0;
      in[760] <= 0;
      in[761] <= 0;
      in[762] <= 0;
      in[763] <= 0;
      in[764] <= 0;
      in[765] <= 0;
      in[766] <= 0;
      in[767] <= 0;
      in[768] <= 0;
      in[769] <= 0;
      in[770] <= 0;
      in[771] <= 0;
      in[772] <= 0;
      in[773] <= 0;
      in[774] <= 0;
      in[775] <= 0;
      in[776] <= 0;
      in[777] <= 0;
      in[778] <= 0;
      in[779] <= 0;
      in[780] <= 0;
      in[781] <= 0;
      in[782] <= 0;
      in[783] <= 0;
      in[784] <= 0;
      in[785] <= 0;
      in[786] <= 0;
      in[787] <= 0;
      in[788] <= 0;
      in[789] <= 0;
      in[790] <= 0;
      in[791] <= 0;
      in[792] <= 0;
      in[793] <= 0;
      in[794] <= 0;
      in[795] <= 0;
      in[796] <= 0;
      in[797] <= 0;
      in[798] <= 0;
      in[799] <= 0;
      in[800] <= 0;
      in[801] <= 0;
      in[802] <= 0;
      in[803] <= 0;
      in[804] <= 0;
      in[805] <= 0;
      in[806] <= 0;
      in[807] <= 0;
      in[808] <= 0;
      in[809] <= 0;
      in[810] <= 0;
      in[811] <= 0;
      in[812] <= 0;
      in[813] <= 0;
      in[814] <= 0;
      in[815] <= 0;
      in[816] <= 0;
      in[817] <= 0;
      in[818] <= 0;
      in[819] <= 0;
      in[820] <= 0;
      in[821] <= 0;
      in[822] <= 0;
      in[823] <= 0;
      in[824] <= 0;
      in[825] <= 0;
      in[826] <= 0;
      in[827] <= 0;
      in[828] <= 0;
      in[829] <= 0;
      in[830] <= 0;
      in[831] <= 0;
      in[832] <= 0;
      in[833] <= 0;
      in[834] <= 0;
      in[835] <= 0;
      in[836] <= 0;
      in[837] <= 0;
      in[838] <= 0;
      in[839] <= 0;
      in[840] <= 0;
      in[841] <= 0;
      in[842] <= 0;
      in[843] <= 0;
      in[844] <= 0;
      in[845] <= 0;
      in[846] <= 0;
      in[847] <= 0;
      in[848] <= 0;
      in[849] <= 0;
      in[850] <= 0;
      in[851] <= 0;
      in[852] <= 0;
      in[853] <= 0;
      in[854] <= 0;
      in[855] <= 0;
      in[856] <= 0;
      in[857] <= 0;
      in[858] <= 0;
      in[859] <= 0;
      in[860] <= 0;
      in[861] <= 0;
      in[862] <= 0;
      in[863] <= 0;
      in[864] <= 0;
      in[865] <= 0;
      in[866] <= 0;
      in[867] <= 0;
      in[868] <= 0;
      in[869] <= 0;
      in[870] <= 0;
      in[871] <= 0;
      in[872] <= 0;
      in[873] <= 0;
      in[874] <= 0;
      in[875] <= 0;
      in[876] <= 0;
      in[877] <= 0;
      in[878] <= 0;
      in[879] <= 0;
      in[880] <= 0;
      in[881] <= 0;
      in[882] <= 0;
      in[883] <= 0;
      in[884] <= 0;
      in[885] <= 0;
      in[886] <= 0;
      in[887] <= 0;
      in[888] <= 0;
      in[889] <= 0;
      in[890] <= 0;
      in[891] <= 0;
      in[892] <= 0;
      in[893] <= 0;
      in[894] <= 0;
      in[895] <= 0;
      in[896] <= 0;
      in[897] <= 0;
      in[898] <= 0;
      in[899] <= 0;
      in[900] <= 0;
      in[901] <= 0;
      in[902] <= 0;
      in[903] <= 0;
      in[904] <= 0;
      in[905] <= 0;
      in[906] <= 0;
      in[907] <= 0;
      in[908] <= 0;
      in[909] <= 0;
      in[910] <= 0;
      in[911] <= 0;
      in[912] <= 0;
      in[913] <= 0;
      in[914] <= 0;
      in[915] <= 0;
      in[916] <= 0;
      in[917] <= 0;
      in[918] <= 0;
      in[919] <= 0;
      in[920] <= 0;
      in[921] <= 0;
      in[922] <= 0;
      in[923] <= 0;
      in[924] <= 0;
      in[925] <= 0;
      in[926] <= 0;
      in[927] <= 0;
      in[928] <= 0;
      in[929] <= 0;
      in[930] <= 0;
      in[931] <= 0;
      in[932] <= 0;
      in[933] <= 0;
      in[934] <= 0;
      in[935] <= 0;
      in[936] <= 0;
      in[937] <= 0;
      in[938] <= 0;
      in[939] <= 0;
      in[940] <= 0;
      in[941] <= 0;
      in[942] <= 0;
      in[943] <= 0;
      in[944] <= 0;
      in[945] <= 0;
      in[946] <= 0;
      in[947] <= 0;
      in[948] <= 0;
      in[949] <= 0;
      in[950] <= 0;
      in[951] <= 0;
      in[952] <= 0;
      in[953] <= 0;
      in[954] <= 0;
      in[955] <= 0;
      in[956] <= 0;
      in[957] <= 0;
      in[958] <= 0;
      in[959] <= 0;
      in[960] <= 0;
      in[961] <= 0;
      in[962] <= 0;
      in[963] <= 0;
      in[964] <= 0;
      in[965] <= 0;
      in[966] <= 0;
      in[967] <= 0;
      in[968] <= 0;
      in[969] <= 0;
      in[970] <= 0;
      in[971] <= 0;
      in[972] <= 0;
      in[973] <= 0;
      in[974] <= 0;
      in[975] <= 0;
      in[976] <= 0;
      in[977] <= 0;
      in[978] <= 0;
      in[979] <= 0;
      in[980] <= 0;
      in[981] <= 0;
      in[982] <= 0;
      in[983] <= 0;
      in[984] <= 0;
      in[985] <= 0;
      in[986] <= 0;
      in[987] <= 0;
      in[988] <= 0;
      in[989] <= 0;
      in[990] <= 0;
      in[991] <= 0;
      in[992] <= 0;
      in[993] <= 0;
      in[994] <= 0;
      in[995] <= 0;
      in[996] <= 0;
      in[997] <= 0;
      in[998] <= 0;
      in[999] <= 0;
      in[1000] <= 0;
      in[1001] <= 0;
      in[1002] <= 0;
      in[1003] <= 0;
      in[1004] <= 0;
      in[1005] <= 0;
      in[1006] <= 0;
      in[1007] <= 0;
      in[1008] <= 0;
      in[1009] <= 0;
      in[1010] <= 0;
      in[1011] <= 0;
      in[1012] <= 0;
      in[1013] <= 0;
      in[1014] <= 0;
      in[1015] <= 0;
      in[1016] <= 0;
      in[1017] <= 0;
      in[1018] <= 0;
      in[1019] <= 0;
      in[1020] <= 0;
      in[1021] <= 0;
      in[1022] <= 0;
      in[1023] <= 0;
      next <= 0;
      reset <= 0;

      @(posedge clk);
      reset <= 1;
      @(posedge clk);
      reset <= 0;
      @(posedge clk);
      @(posedge clk);
      // Wait until next_out goes high, then wait one clock cycle and begin receiving data
      @(posedge next_out);
      @(posedge clk); #1;
      $display("--- begin output 1---");

      for (m=0; m < 0; m=m+1) begin
         $display("%x", Y0);
         $display("%x", Y1);
         $display("%x", Y2);
         $display("%x", Y3);
         $display("%x", Y4);
         $display("%x", Y5);
         $display("%x", Y6);
         $display("%x", Y7);
         $display("%x", Y8);
         $display("%x", Y9);
         $display("%x", Y10);
         $display("%x", Y11);
         $display("%x", Y12);
         $display("%x", Y13);
         $display("%x", Y14);
         $display("%x", Y15);
         $display("%x", Y16);
         $display("%x", Y17);
         $display("%x", Y18);
         $display("%x", Y19);
         $display("%x", Y20);
         $display("%x", Y21);
         $display("%x", Y22);
         $display("%x", Y23);
         $display("%x", Y24);
         $display("%x", Y25);
         $display("%x", Y26);
         $display("%x", Y27);
         $display("%x", Y28);
         $display("%x", Y29);
         $display("%x", Y30);
         $display("%x", Y31);
         $display("%x", Y32);
         $display("%x", Y33);
         $display("%x", Y34);
         $display("%x", Y35);
         $display("%x", Y36);
         $display("%x", Y37);
         $display("%x", Y38);
         $display("%x", Y39);
         $display("%x", Y40);
         $display("%x", Y41);
         $display("%x", Y42);
         $display("%x", Y43);
         $display("%x", Y44);
         $display("%x", Y45);
         $display("%x", Y46);
         $display("%x", Y47);
         $display("%x", Y48);
         $display("%x", Y49);
         $display("%x", Y50);
         $display("%x", Y51);
         $display("%x", Y52);
         $display("%x", Y53);
         $display("%x", Y54);
         $display("%x", Y55);
         $display("%x", Y56);
         $display("%x", Y57);
         $display("%x", Y58);
         $display("%x", Y59);
         $display("%x", Y60);
         $display("%x", Y61);
         $display("%x", Y62);
         $display("%x", Y63);
         $display("%x", Y64);
         $display("%x", Y65);
         $display("%x", Y66);
         $display("%x", Y67);
         $display("%x", Y68);
         $display("%x", Y69);
         $display("%x", Y70);
         $display("%x", Y71);
         $display("%x", Y72);
         $display("%x", Y73);
         $display("%x", Y74);
         $display("%x", Y75);
         $display("%x", Y76);
         $display("%x", Y77);
         $display("%x", Y78);
         $display("%x", Y79);
         $display("%x", Y80);
         $display("%x", Y81);
         $display("%x", Y82);
         $display("%x", Y83);
         $display("%x", Y84);
         $display("%x", Y85);
         $display("%x", Y86);
         $display("%x", Y87);
         $display("%x", Y88);
         $display("%x", Y89);
         $display("%x", Y90);
         $display("%x", Y91);
         $display("%x", Y92);
         $display("%x", Y93);
         $display("%x", Y94);
         $display("%x", Y95);
         $display("%x", Y96);
         $display("%x", Y97);
         $display("%x", Y98);
         $display("%x", Y99);
         $display("%x", Y100);
         $display("%x", Y101);
         $display("%x", Y102);
         $display("%x", Y103);
         $display("%x", Y104);
         $display("%x", Y105);
         $display("%x", Y106);
         $display("%x", Y107);
         $display("%x", Y108);
         $display("%x", Y109);
         $display("%x", Y110);
         $display("%x", Y111);
         $display("%x", Y112);
         $display("%x", Y113);
         $display("%x", Y114);
         $display("%x", Y115);
         $display("%x", Y116);
         $display("%x", Y117);
         $display("%x", Y118);
         $display("%x", Y119);
         $display("%x", Y120);
         $display("%x", Y121);
         $display("%x", Y122);
         $display("%x", Y123);
         $display("%x", Y124);
         $display("%x", Y125);
         $display("%x", Y126);
         $display("%x", Y127);
         $display("%x", Y128);
         $display("%x", Y129);
         $display("%x", Y130);
         $display("%x", Y131);
         $display("%x", Y132);
         $display("%x", Y133);
         $display("%x", Y134);
         $display("%x", Y135);
         $display("%x", Y136);
         $display("%x", Y137);
         $display("%x", Y138);
         $display("%x", Y139);
         $display("%x", Y140);
         $display("%x", Y141);
         $display("%x", Y142);
         $display("%x", Y143);
         $display("%x", Y144);
         $display("%x", Y145);
         $display("%x", Y146);
         $display("%x", Y147);
         $display("%x", Y148);
         $display("%x", Y149);
         $display("%x", Y150);
         $display("%x", Y151);
         $display("%x", Y152);
         $display("%x", Y153);
         $display("%x", Y154);
         $display("%x", Y155);
         $display("%x", Y156);
         $display("%x", Y157);
         $display("%x", Y158);
         $display("%x", Y159);
         $display("%x", Y160);
         $display("%x", Y161);
         $display("%x", Y162);
         $display("%x", Y163);
         $display("%x", Y164);
         $display("%x", Y165);
         $display("%x", Y166);
         $display("%x", Y167);
         $display("%x", Y168);
         $display("%x", Y169);
         $display("%x", Y170);
         $display("%x", Y171);
         $display("%x", Y172);
         $display("%x", Y173);
         $display("%x", Y174);
         $display("%x", Y175);
         $display("%x", Y176);
         $display("%x", Y177);
         $display("%x", Y178);
         $display("%x", Y179);
         $display("%x", Y180);
         $display("%x", Y181);
         $display("%x", Y182);
         $display("%x", Y183);
         $display("%x", Y184);
         $display("%x", Y185);
         $display("%x", Y186);
         $display("%x", Y187);
         $display("%x", Y188);
         $display("%x", Y189);
         $display("%x", Y190);
         $display("%x", Y191);
         $display("%x", Y192);
         $display("%x", Y193);
         $display("%x", Y194);
         $display("%x", Y195);
         $display("%x", Y196);
         $display("%x", Y197);
         $display("%x", Y198);
         $display("%x", Y199);
         $display("%x", Y200);
         $display("%x", Y201);
         $display("%x", Y202);
         $display("%x", Y203);
         $display("%x", Y204);
         $display("%x", Y205);
         $display("%x", Y206);
         $display("%x", Y207);
         $display("%x", Y208);
         $display("%x", Y209);
         $display("%x", Y210);
         $display("%x", Y211);
         $display("%x", Y212);
         $display("%x", Y213);
         $display("%x", Y214);
         $display("%x", Y215);
         $display("%x", Y216);
         $display("%x", Y217);
         $display("%x", Y218);
         $display("%x", Y219);
         $display("%x", Y220);
         $display("%x", Y221);
         $display("%x", Y222);
         $display("%x", Y223);
         $display("%x", Y224);
         $display("%x", Y225);
         $display("%x", Y226);
         $display("%x", Y227);
         $display("%x", Y228);
         $display("%x", Y229);
         $display("%x", Y230);
         $display("%x", Y231);
         $display("%x", Y232);
         $display("%x", Y233);
         $display("%x", Y234);
         $display("%x", Y235);
         $display("%x", Y236);
         $display("%x", Y237);
         $display("%x", Y238);
         $display("%x", Y239);
         $display("%x", Y240);
         $display("%x", Y241);
         $display("%x", Y242);
         $display("%x", Y243);
         $display("%x", Y244);
         $display("%x", Y245);
         $display("%x", Y246);
         $display("%x", Y247);
         $display("%x", Y248);
         $display("%x", Y249);
         $display("%x", Y250);
         $display("%x", Y251);
         $display("%x", Y252);
         $display("%x", Y253);
         $display("%x", Y254);
         $display("%x", Y255);
         $display("%x", Y256);
         $display("%x", Y257);
         $display("%x", Y258);
         $display("%x", Y259);
         $display("%x", Y260);
         $display("%x", Y261);
         $display("%x", Y262);
         $display("%x", Y263);
         $display("%x", Y264);
         $display("%x", Y265);
         $display("%x", Y266);
         $display("%x", Y267);
         $display("%x", Y268);
         $display("%x", Y269);
         $display("%x", Y270);
         $display("%x", Y271);
         $display("%x", Y272);
         $display("%x", Y273);
         $display("%x", Y274);
         $display("%x", Y275);
         $display("%x", Y276);
         $display("%x", Y277);
         $display("%x", Y278);
         $display("%x", Y279);
         $display("%x", Y280);
         $display("%x", Y281);
         $display("%x", Y282);
         $display("%x", Y283);
         $display("%x", Y284);
         $display("%x", Y285);
         $display("%x", Y286);
         $display("%x", Y287);
         $display("%x", Y288);
         $display("%x", Y289);
         $display("%x", Y290);
         $display("%x", Y291);
         $display("%x", Y292);
         $display("%x", Y293);
         $display("%x", Y294);
         $display("%x", Y295);
         $display("%x", Y296);
         $display("%x", Y297);
         $display("%x", Y298);
         $display("%x", Y299);
         $display("%x", Y300);
         $display("%x", Y301);
         $display("%x", Y302);
         $display("%x", Y303);
         $display("%x", Y304);
         $display("%x", Y305);
         $display("%x", Y306);
         $display("%x", Y307);
         $display("%x", Y308);
         $display("%x", Y309);
         $display("%x", Y310);
         $display("%x", Y311);
         $display("%x", Y312);
         $display("%x", Y313);
         $display("%x", Y314);
         $display("%x", Y315);
         $display("%x", Y316);
         $display("%x", Y317);
         $display("%x", Y318);
         $display("%x", Y319);
         $display("%x", Y320);
         $display("%x", Y321);
         $display("%x", Y322);
         $display("%x", Y323);
         $display("%x", Y324);
         $display("%x", Y325);
         $display("%x", Y326);
         $display("%x", Y327);
         $display("%x", Y328);
         $display("%x", Y329);
         $display("%x", Y330);
         $display("%x", Y331);
         $display("%x", Y332);
         $display("%x", Y333);
         $display("%x", Y334);
         $display("%x", Y335);
         $display("%x", Y336);
         $display("%x", Y337);
         $display("%x", Y338);
         $display("%x", Y339);
         $display("%x", Y340);
         $display("%x", Y341);
         $display("%x", Y342);
         $display("%x", Y343);
         $display("%x", Y344);
         $display("%x", Y345);
         $display("%x", Y346);
         $display("%x", Y347);
         $display("%x", Y348);
         $display("%x", Y349);
         $display("%x", Y350);
         $display("%x", Y351);
         $display("%x", Y352);
         $display("%x", Y353);
         $display("%x", Y354);
         $display("%x", Y355);
         $display("%x", Y356);
         $display("%x", Y357);
         $display("%x", Y358);
         $display("%x", Y359);
         $display("%x", Y360);
         $display("%x", Y361);
         $display("%x", Y362);
         $display("%x", Y363);
         $display("%x", Y364);
         $display("%x", Y365);
         $display("%x", Y366);
         $display("%x", Y367);
         $display("%x", Y368);
         $display("%x", Y369);
         $display("%x", Y370);
         $display("%x", Y371);
         $display("%x", Y372);
         $display("%x", Y373);
         $display("%x", Y374);
         $display("%x", Y375);
         $display("%x", Y376);
         $display("%x", Y377);
         $display("%x", Y378);
         $display("%x", Y379);
         $display("%x", Y380);
         $display("%x", Y381);
         $display("%x", Y382);
         $display("%x", Y383);
         $display("%x", Y384);
         $display("%x", Y385);
         $display("%x", Y386);
         $display("%x", Y387);
         $display("%x", Y388);
         $display("%x", Y389);
         $display("%x", Y390);
         $display("%x", Y391);
         $display("%x", Y392);
         $display("%x", Y393);
         $display("%x", Y394);
         $display("%x", Y395);
         $display("%x", Y396);
         $display("%x", Y397);
         $display("%x", Y398);
         $display("%x", Y399);
         $display("%x", Y400);
         $display("%x", Y401);
         $display("%x", Y402);
         $display("%x", Y403);
         $display("%x", Y404);
         $display("%x", Y405);
         $display("%x", Y406);
         $display("%x", Y407);
         $display("%x", Y408);
         $display("%x", Y409);
         $display("%x", Y410);
         $display("%x", Y411);
         $display("%x", Y412);
         $display("%x", Y413);
         $display("%x", Y414);
         $display("%x", Y415);
         $display("%x", Y416);
         $display("%x", Y417);
         $display("%x", Y418);
         $display("%x", Y419);
         $display("%x", Y420);
         $display("%x", Y421);
         $display("%x", Y422);
         $display("%x", Y423);
         $display("%x", Y424);
         $display("%x", Y425);
         $display("%x", Y426);
         $display("%x", Y427);
         $display("%x", Y428);
         $display("%x", Y429);
         $display("%x", Y430);
         $display("%x", Y431);
         $display("%x", Y432);
         $display("%x", Y433);
         $display("%x", Y434);
         $display("%x", Y435);
         $display("%x", Y436);
         $display("%x", Y437);
         $display("%x", Y438);
         $display("%x", Y439);
         $display("%x", Y440);
         $display("%x", Y441);
         $display("%x", Y442);
         $display("%x", Y443);
         $display("%x", Y444);
         $display("%x", Y445);
         $display("%x", Y446);
         $display("%x", Y447);
         $display("%x", Y448);
         $display("%x", Y449);
         $display("%x", Y450);
         $display("%x", Y451);
         $display("%x", Y452);
         $display("%x", Y453);
         $display("%x", Y454);
         $display("%x", Y455);
         $display("%x", Y456);
         $display("%x", Y457);
         $display("%x", Y458);
         $display("%x", Y459);
         $display("%x", Y460);
         $display("%x", Y461);
         $display("%x", Y462);
         $display("%x", Y463);
         $display("%x", Y464);
         $display("%x", Y465);
         $display("%x", Y466);
         $display("%x", Y467);
         $display("%x", Y468);
         $display("%x", Y469);
         $display("%x", Y470);
         $display("%x", Y471);
         $display("%x", Y472);
         $display("%x", Y473);
         $display("%x", Y474);
         $display("%x", Y475);
         $display("%x", Y476);
         $display("%x", Y477);
         $display("%x", Y478);
         $display("%x", Y479);
         $display("%x", Y480);
         $display("%x", Y481);
         $display("%x", Y482);
         $display("%x", Y483);
         $display("%x", Y484);
         $display("%x", Y485);
         $display("%x", Y486);
         $display("%x", Y487);
         $display("%x", Y488);
         $display("%x", Y489);
         $display("%x", Y490);
         $display("%x", Y491);
         $display("%x", Y492);
         $display("%x", Y493);
         $display("%x", Y494);
         $display("%x", Y495);
         $display("%x", Y496);
         $display("%x", Y497);
         $display("%x", Y498);
         $display("%x", Y499);
         $display("%x", Y500);
         $display("%x", Y501);
         $display("%x", Y502);
         $display("%x", Y503);
         $display("%x", Y504);
         $display("%x", Y505);
         $display("%x", Y506);
         $display("%x", Y507);
         $display("%x", Y508);
         $display("%x", Y509);
         $display("%x", Y510);
         $display("%x", Y511);
         $display("%x", Y512);
         $display("%x", Y513);
         $display("%x", Y514);
         $display("%x", Y515);
         $display("%x", Y516);
         $display("%x", Y517);
         $display("%x", Y518);
         $display("%x", Y519);
         $display("%x", Y520);
         $display("%x", Y521);
         $display("%x", Y522);
         $display("%x", Y523);
         $display("%x", Y524);
         $display("%x", Y525);
         $display("%x", Y526);
         $display("%x", Y527);
         $display("%x", Y528);
         $display("%x", Y529);
         $display("%x", Y530);
         $display("%x", Y531);
         $display("%x", Y532);
         $display("%x", Y533);
         $display("%x", Y534);
         $display("%x", Y535);
         $display("%x", Y536);
         $display("%x", Y537);
         $display("%x", Y538);
         $display("%x", Y539);
         $display("%x", Y540);
         $display("%x", Y541);
         $display("%x", Y542);
         $display("%x", Y543);
         $display("%x", Y544);
         $display("%x", Y545);
         $display("%x", Y546);
         $display("%x", Y547);
         $display("%x", Y548);
         $display("%x", Y549);
         $display("%x", Y550);
         $display("%x", Y551);
         $display("%x", Y552);
         $display("%x", Y553);
         $display("%x", Y554);
         $display("%x", Y555);
         $display("%x", Y556);
         $display("%x", Y557);
         $display("%x", Y558);
         $display("%x", Y559);
         $display("%x", Y560);
         $display("%x", Y561);
         $display("%x", Y562);
         $display("%x", Y563);
         $display("%x", Y564);
         $display("%x", Y565);
         $display("%x", Y566);
         $display("%x", Y567);
         $display("%x", Y568);
         $display("%x", Y569);
         $display("%x", Y570);
         $display("%x", Y571);
         $display("%x", Y572);
         $display("%x", Y573);
         $display("%x", Y574);
         $display("%x", Y575);
         $display("%x", Y576);
         $display("%x", Y577);
         $display("%x", Y578);
         $display("%x", Y579);
         $display("%x", Y580);
         $display("%x", Y581);
         $display("%x", Y582);
         $display("%x", Y583);
         $display("%x", Y584);
         $display("%x", Y585);
         $display("%x", Y586);
         $display("%x", Y587);
         $display("%x", Y588);
         $display("%x", Y589);
         $display("%x", Y590);
         $display("%x", Y591);
         $display("%x", Y592);
         $display("%x", Y593);
         $display("%x", Y594);
         $display("%x", Y595);
         $display("%x", Y596);
         $display("%x", Y597);
         $display("%x", Y598);
         $display("%x", Y599);
         $display("%x", Y600);
         $display("%x", Y601);
         $display("%x", Y602);
         $display("%x", Y603);
         $display("%x", Y604);
         $display("%x", Y605);
         $display("%x", Y606);
         $display("%x", Y607);
         $display("%x", Y608);
         $display("%x", Y609);
         $display("%x", Y610);
         $display("%x", Y611);
         $display("%x", Y612);
         $display("%x", Y613);
         $display("%x", Y614);
         $display("%x", Y615);
         $display("%x", Y616);
         $display("%x", Y617);
         $display("%x", Y618);
         $display("%x", Y619);
         $display("%x", Y620);
         $display("%x", Y621);
         $display("%x", Y622);
         $display("%x", Y623);
         $display("%x", Y624);
         $display("%x", Y625);
         $display("%x", Y626);
         $display("%x", Y627);
         $display("%x", Y628);
         $display("%x", Y629);
         $display("%x", Y630);
         $display("%x", Y631);
         $display("%x", Y632);
         $display("%x", Y633);
         $display("%x", Y634);
         $display("%x", Y635);
         $display("%x", Y636);
         $display("%x", Y637);
         $display("%x", Y638);
         $display("%x", Y639);
         $display("%x", Y640);
         $display("%x", Y641);
         $display("%x", Y642);
         $display("%x", Y643);
         $display("%x", Y644);
         $display("%x", Y645);
         $display("%x", Y646);
         $display("%x", Y647);
         $display("%x", Y648);
         $display("%x", Y649);
         $display("%x", Y650);
         $display("%x", Y651);
         $display("%x", Y652);
         $display("%x", Y653);
         $display("%x", Y654);
         $display("%x", Y655);
         $display("%x", Y656);
         $display("%x", Y657);
         $display("%x", Y658);
         $display("%x", Y659);
         $display("%x", Y660);
         $display("%x", Y661);
         $display("%x", Y662);
         $display("%x", Y663);
         $display("%x", Y664);
         $display("%x", Y665);
         $display("%x", Y666);
         $display("%x", Y667);
         $display("%x", Y668);
         $display("%x", Y669);
         $display("%x", Y670);
         $display("%x", Y671);
         $display("%x", Y672);
         $display("%x", Y673);
         $display("%x", Y674);
         $display("%x", Y675);
         $display("%x", Y676);
         $display("%x", Y677);
         $display("%x", Y678);
         $display("%x", Y679);
         $display("%x", Y680);
         $display("%x", Y681);
         $display("%x", Y682);
         $display("%x", Y683);
         $display("%x", Y684);
         $display("%x", Y685);
         $display("%x", Y686);
         $display("%x", Y687);
         $display("%x", Y688);
         $display("%x", Y689);
         $display("%x", Y690);
         $display("%x", Y691);
         $display("%x", Y692);
         $display("%x", Y693);
         $display("%x", Y694);
         $display("%x", Y695);
         $display("%x", Y696);
         $display("%x", Y697);
         $display("%x", Y698);
         $display("%x", Y699);
         $display("%x", Y700);
         $display("%x", Y701);
         $display("%x", Y702);
         $display("%x", Y703);
         $display("%x", Y704);
         $display("%x", Y705);
         $display("%x", Y706);
         $display("%x", Y707);
         $display("%x", Y708);
         $display("%x", Y709);
         $display("%x", Y710);
         $display("%x", Y711);
         $display("%x", Y712);
         $display("%x", Y713);
         $display("%x", Y714);
         $display("%x", Y715);
         $display("%x", Y716);
         $display("%x", Y717);
         $display("%x", Y718);
         $display("%x", Y719);
         $display("%x", Y720);
         $display("%x", Y721);
         $display("%x", Y722);
         $display("%x", Y723);
         $display("%x", Y724);
         $display("%x", Y725);
         $display("%x", Y726);
         $display("%x", Y727);
         $display("%x", Y728);
         $display("%x", Y729);
         $display("%x", Y730);
         $display("%x", Y731);
         $display("%x", Y732);
         $display("%x", Y733);
         $display("%x", Y734);
         $display("%x", Y735);
         $display("%x", Y736);
         $display("%x", Y737);
         $display("%x", Y738);
         $display("%x", Y739);
         $display("%x", Y740);
         $display("%x", Y741);
         $display("%x", Y742);
         $display("%x", Y743);
         $display("%x", Y744);
         $display("%x", Y745);
         $display("%x", Y746);
         $display("%x", Y747);
         $display("%x", Y748);
         $display("%x", Y749);
         $display("%x", Y750);
         $display("%x", Y751);
         $display("%x", Y752);
         $display("%x", Y753);
         $display("%x", Y754);
         $display("%x", Y755);
         $display("%x", Y756);
         $display("%x", Y757);
         $display("%x", Y758);
         $display("%x", Y759);
         $display("%x", Y760);
         $display("%x", Y761);
         $display("%x", Y762);
         $display("%x", Y763);
         $display("%x", Y764);
         $display("%x", Y765);
         $display("%x", Y766);
         $display("%x", Y767);
         $display("%x", Y768);
         $display("%x", Y769);
         $display("%x", Y770);
         $display("%x", Y771);
         $display("%x", Y772);
         $display("%x", Y773);
         $display("%x", Y774);
         $display("%x", Y775);
         $display("%x", Y776);
         $display("%x", Y777);
         $display("%x", Y778);
         $display("%x", Y779);
         $display("%x", Y780);
         $display("%x", Y781);
         $display("%x", Y782);
         $display("%x", Y783);
         $display("%x", Y784);
         $display("%x", Y785);
         $display("%x", Y786);
         $display("%x", Y787);
         $display("%x", Y788);
         $display("%x", Y789);
         $display("%x", Y790);
         $display("%x", Y791);
         $display("%x", Y792);
         $display("%x", Y793);
         $display("%x", Y794);
         $display("%x", Y795);
         $display("%x", Y796);
         $display("%x", Y797);
         $display("%x", Y798);
         $display("%x", Y799);
         $display("%x", Y800);
         $display("%x", Y801);
         $display("%x", Y802);
         $display("%x", Y803);
         $display("%x", Y804);
         $display("%x", Y805);
         $display("%x", Y806);
         $display("%x", Y807);
         $display("%x", Y808);
         $display("%x", Y809);
         $display("%x", Y810);
         $display("%x", Y811);
         $display("%x", Y812);
         $display("%x", Y813);
         $display("%x", Y814);
         $display("%x", Y815);
         $display("%x", Y816);
         $display("%x", Y817);
         $display("%x", Y818);
         $display("%x", Y819);
         $display("%x", Y820);
         $display("%x", Y821);
         $display("%x", Y822);
         $display("%x", Y823);
         $display("%x", Y824);
         $display("%x", Y825);
         $display("%x", Y826);
         $display("%x", Y827);
         $display("%x", Y828);
         $display("%x", Y829);
         $display("%x", Y830);
         $display("%x", Y831);
         $display("%x", Y832);
         $display("%x", Y833);
         $display("%x", Y834);
         $display("%x", Y835);
         $display("%x", Y836);
         $display("%x", Y837);
         $display("%x", Y838);
         $display("%x", Y839);
         $display("%x", Y840);
         $display("%x", Y841);
         $display("%x", Y842);
         $display("%x", Y843);
         $display("%x", Y844);
         $display("%x", Y845);
         $display("%x", Y846);
         $display("%x", Y847);
         $display("%x", Y848);
         $display("%x", Y849);
         $display("%x", Y850);
         $display("%x", Y851);
         $display("%x", Y852);
         $display("%x", Y853);
         $display("%x", Y854);
         $display("%x", Y855);
         $display("%x", Y856);
         $display("%x", Y857);
         $display("%x", Y858);
         $display("%x", Y859);
         $display("%x", Y860);
         $display("%x", Y861);
         $display("%x", Y862);
         $display("%x", Y863);
         $display("%x", Y864);
         $display("%x", Y865);
         $display("%x", Y866);
         $display("%x", Y867);
         $display("%x", Y868);
         $display("%x", Y869);
         $display("%x", Y870);
         $display("%x", Y871);
         $display("%x", Y872);
         $display("%x", Y873);
         $display("%x", Y874);
         $display("%x", Y875);
         $display("%x", Y876);
         $display("%x", Y877);
         $display("%x", Y878);
         $display("%x", Y879);
         $display("%x", Y880);
         $display("%x", Y881);
         $display("%x", Y882);
         $display("%x", Y883);
         $display("%x", Y884);
         $display("%x", Y885);
         $display("%x", Y886);
         $display("%x", Y887);
         $display("%x", Y888);
         $display("%x", Y889);
         $display("%x", Y890);
         $display("%x", Y891);
         $display("%x", Y892);
         $display("%x", Y893);
         $display("%x", Y894);
         $display("%x", Y895);
         $display("%x", Y896);
         $display("%x", Y897);
         $display("%x", Y898);
         $display("%x", Y899);
         $display("%x", Y900);
         $display("%x", Y901);
         $display("%x", Y902);
         $display("%x", Y903);
         $display("%x", Y904);
         $display("%x", Y905);
         $display("%x", Y906);
         $display("%x", Y907);
         $display("%x", Y908);
         $display("%x", Y909);
         $display("%x", Y910);
         $display("%x", Y911);
         $display("%x", Y912);
         $display("%x", Y913);
         $display("%x", Y914);
         $display("%x", Y915);
         $display("%x", Y916);
         $display("%x", Y917);
         $display("%x", Y918);
         $display("%x", Y919);
         $display("%x", Y920);
         $display("%x", Y921);
         $display("%x", Y922);
         $display("%x", Y923);
         $display("%x", Y924);
         $display("%x", Y925);
         $display("%x", Y926);
         $display("%x", Y927);
         $display("%x", Y928);
         $display("%x", Y929);
         $display("%x", Y930);
         $display("%x", Y931);
         $display("%x", Y932);
         $display("%x", Y933);
         $display("%x", Y934);
         $display("%x", Y935);
         $display("%x", Y936);
         $display("%x", Y937);
         $display("%x", Y938);
         $display("%x", Y939);
         $display("%x", Y940);
         $display("%x", Y941);
         $display("%x", Y942);
         $display("%x", Y943);
         $display("%x", Y944);
         $display("%x", Y945);
         $display("%x", Y946);
         $display("%x", Y947);
         $display("%x", Y948);
         $display("%x", Y949);
         $display("%x", Y950);
         $display("%x", Y951);
         $display("%x", Y952);
         $display("%x", Y953);
         $display("%x", Y954);
         $display("%x", Y955);
         $display("%x", Y956);
         $display("%x", Y957);
         $display("%x", Y958);
         $display("%x", Y959);
         $display("%x", Y960);
         $display("%x", Y961);
         $display("%x", Y962);
         $display("%x", Y963);
         $display("%x", Y964);
         $display("%x", Y965);
         $display("%x", Y966);
         $display("%x", Y967);
         $display("%x", Y968);
         $display("%x", Y969);
         $display("%x", Y970);
         $display("%x", Y971);
         $display("%x", Y972);
         $display("%x", Y973);
         $display("%x", Y974);
         $display("%x", Y975);
         $display("%x", Y976);
         $display("%x", Y977);
         $display("%x", Y978);
         $display("%x", Y979);
         $display("%x", Y980);
         $display("%x", Y981);
         $display("%x", Y982);
         $display("%x", Y983);
         $display("%x", Y984);
         $display("%x", Y985);
         $display("%x", Y986);
         $display("%x", Y987);
         $display("%x", Y988);
         $display("%x", Y989);
         $display("%x", Y990);
         $display("%x", Y991);
         $display("%x", Y992);
         $display("%x", Y993);
         $display("%x", Y994);
         $display("%x", Y995);
         $display("%x", Y996);
         $display("%x", Y997);
         $display("%x", Y998);
         $display("%x", Y999);
         $display("%x", Y1000);
         $display("%x", Y1001);
         $display("%x", Y1002);
         $display("%x", Y1003);
         $display("%x", Y1004);
         $display("%x", Y1005);
         $display("%x", Y1006);
         $display("%x", Y1007);
         $display("%x", Y1008);
         $display("%x", Y1009);
         $display("%x", Y1010);
         $display("%x", Y1011);
         $display("%x", Y1012);
         $display("%x", Y1013);
         $display("%x", Y1014);
         $display("%x", Y1015);
         $display("%x", Y1016);
         $display("%x", Y1017);
         $display("%x", Y1018);
         $display("%x", Y1019);
         $display("%x", Y1020);
         $display("%x", Y1021);
         $display("%x", Y1022);
         $display("%x", Y1023);
         @(posedge clk); #1;
      end
      $display("%x", Y0);
      $display("%x", Y1);
      $display("%x", Y2);
      $display("%x", Y3);
      $display("%x", Y4);
      $display("%x", Y5);
      $display("%x", Y6);
      $display("%x", Y7);
      $display("%x", Y8);
      $display("%x", Y9);
      $display("%x", Y10);
      $display("%x", Y11);
      $display("%x", Y12);
      $display("%x", Y13);
      $display("%x", Y14);
      $display("%x", Y15);
      $display("%x", Y16);
      $display("%x", Y17);
      $display("%x", Y18);
      $display("%x", Y19);
      $display("%x", Y20);
      $display("%x", Y21);
      $display("%x", Y22);
      $display("%x", Y23);
      $display("%x", Y24);
      $display("%x", Y25);
      $display("%x", Y26);
      $display("%x", Y27);
      $display("%x", Y28);
      $display("%x", Y29);
      $display("%x", Y30);
      $display("%x", Y31);
      $display("%x", Y32);
      $display("%x", Y33);
      $display("%x", Y34);
      $display("%x", Y35);
      $display("%x", Y36);
      $display("%x", Y37);
      $display("%x", Y38);
      $display("%x", Y39);
      $display("%x", Y40);
      $display("%x", Y41);
      $display("%x", Y42);
      $display("%x", Y43);
      $display("%x", Y44);
      $display("%x", Y45);
      $display("%x", Y46);
      $display("%x", Y47);
      $display("%x", Y48);
      $display("%x", Y49);
      $display("%x", Y50);
      $display("%x", Y51);
      $display("%x", Y52);
      $display("%x", Y53);
      $display("%x", Y54);
      $display("%x", Y55);
      $display("%x", Y56);
      $display("%x", Y57);
      $display("%x", Y58);
      $display("%x", Y59);
      $display("%x", Y60);
      $display("%x", Y61);
      $display("%x", Y62);
      $display("%x", Y63);
      $display("%x", Y64);
      $display("%x", Y65);
      $display("%x", Y66);
      $display("%x", Y67);
      $display("%x", Y68);
      $display("%x", Y69);
      $display("%x", Y70);
      $display("%x", Y71);
      $display("%x", Y72);
      $display("%x", Y73);
      $display("%x", Y74);
      $display("%x", Y75);
      $display("%x", Y76);
      $display("%x", Y77);
      $display("%x", Y78);
      $display("%x", Y79);
      $display("%x", Y80);
      $display("%x", Y81);
      $display("%x", Y82);
      $display("%x", Y83);
      $display("%x", Y84);
      $display("%x", Y85);
      $display("%x", Y86);
      $display("%x", Y87);
      $display("%x", Y88);
      $display("%x", Y89);
      $display("%x", Y90);
      $display("%x", Y91);
      $display("%x", Y92);
      $display("%x", Y93);
      $display("%x", Y94);
      $display("%x", Y95);
      $display("%x", Y96);
      $display("%x", Y97);
      $display("%x", Y98);
      $display("%x", Y99);
      $display("%x", Y100);
      $display("%x", Y101);
      $display("%x", Y102);
      $display("%x", Y103);
      $display("%x", Y104);
      $display("%x", Y105);
      $display("%x", Y106);
      $display("%x", Y107);
      $display("%x", Y108);
      $display("%x", Y109);
      $display("%x", Y110);
      $display("%x", Y111);
      $display("%x", Y112);
      $display("%x", Y113);
      $display("%x", Y114);
      $display("%x", Y115);
      $display("%x", Y116);
      $display("%x", Y117);
      $display("%x", Y118);
      $display("%x", Y119);
      $display("%x", Y120);
      $display("%x", Y121);
      $display("%x", Y122);
      $display("%x", Y123);
      $display("%x", Y124);
      $display("%x", Y125);
      $display("%x", Y126);
      $display("%x", Y127);
      $display("%x", Y128);
      $display("%x", Y129);
      $display("%x", Y130);
      $display("%x", Y131);
      $display("%x", Y132);
      $display("%x", Y133);
      $display("%x", Y134);
      $display("%x", Y135);
      $display("%x", Y136);
      $display("%x", Y137);
      $display("%x", Y138);
      $display("%x", Y139);
      $display("%x", Y140);
      $display("%x", Y141);
      $display("%x", Y142);
      $display("%x", Y143);
      $display("%x", Y144);
      $display("%x", Y145);
      $display("%x", Y146);
      $display("%x", Y147);
      $display("%x", Y148);
      $display("%x", Y149);
      $display("%x", Y150);
      $display("%x", Y151);
      $display("%x", Y152);
      $display("%x", Y153);
      $display("%x", Y154);
      $display("%x", Y155);
      $display("%x", Y156);
      $display("%x", Y157);
      $display("%x", Y158);
      $display("%x", Y159);
      $display("%x", Y160);
      $display("%x", Y161);
      $display("%x", Y162);
      $display("%x", Y163);
      $display("%x", Y164);
      $display("%x", Y165);
      $display("%x", Y166);
      $display("%x", Y167);
      $display("%x", Y168);
      $display("%x", Y169);
      $display("%x", Y170);
      $display("%x", Y171);
      $display("%x", Y172);
      $display("%x", Y173);
      $display("%x", Y174);
      $display("%x", Y175);
      $display("%x", Y176);
      $display("%x", Y177);
      $display("%x", Y178);
      $display("%x", Y179);
      $display("%x", Y180);
      $display("%x", Y181);
      $display("%x", Y182);
      $display("%x", Y183);
      $display("%x", Y184);
      $display("%x", Y185);
      $display("%x", Y186);
      $display("%x", Y187);
      $display("%x", Y188);
      $display("%x", Y189);
      $display("%x", Y190);
      $display("%x", Y191);
      $display("%x", Y192);
      $display("%x", Y193);
      $display("%x", Y194);
      $display("%x", Y195);
      $display("%x", Y196);
      $display("%x", Y197);
      $display("%x", Y198);
      $display("%x", Y199);
      $display("%x", Y200);
      $display("%x", Y201);
      $display("%x", Y202);
      $display("%x", Y203);
      $display("%x", Y204);
      $display("%x", Y205);
      $display("%x", Y206);
      $display("%x", Y207);
      $display("%x", Y208);
      $display("%x", Y209);
      $display("%x", Y210);
      $display("%x", Y211);
      $display("%x", Y212);
      $display("%x", Y213);
      $display("%x", Y214);
      $display("%x", Y215);
      $display("%x", Y216);
      $display("%x", Y217);
      $display("%x", Y218);
      $display("%x", Y219);
      $display("%x", Y220);
      $display("%x", Y221);
      $display("%x", Y222);
      $display("%x", Y223);
      $display("%x", Y224);
      $display("%x", Y225);
      $display("%x", Y226);
      $display("%x", Y227);
      $display("%x", Y228);
      $display("%x", Y229);
      $display("%x", Y230);
      $display("%x", Y231);
      $display("%x", Y232);
      $display("%x", Y233);
      $display("%x", Y234);
      $display("%x", Y235);
      $display("%x", Y236);
      $display("%x", Y237);
      $display("%x", Y238);
      $display("%x", Y239);
      $display("%x", Y240);
      $display("%x", Y241);
      $display("%x", Y242);
      $display("%x", Y243);
      $display("%x", Y244);
      $display("%x", Y245);
      $display("%x", Y246);
      $display("%x", Y247);
      $display("%x", Y248);
      $display("%x", Y249);
      $display("%x", Y250);
      $display("%x", Y251);
      $display("%x", Y252);
      $display("%x", Y253);
      $display("%x", Y254);
      $display("%x", Y255);
      $display("%x", Y256);
      $display("%x", Y257);
      $display("%x", Y258);
      $display("%x", Y259);
      $display("%x", Y260);
      $display("%x", Y261);
      $display("%x", Y262);
      $display("%x", Y263);
      $display("%x", Y264);
      $display("%x", Y265);
      $display("%x", Y266);
      $display("%x", Y267);
      $display("%x", Y268);
      $display("%x", Y269);
      $display("%x", Y270);
      $display("%x", Y271);
      $display("%x", Y272);
      $display("%x", Y273);
      $display("%x", Y274);
      $display("%x", Y275);
      $display("%x", Y276);
      $display("%x", Y277);
      $display("%x", Y278);
      $display("%x", Y279);
      $display("%x", Y280);
      $display("%x", Y281);
      $display("%x", Y282);
      $display("%x", Y283);
      $display("%x", Y284);
      $display("%x", Y285);
      $display("%x", Y286);
      $display("%x", Y287);
      $display("%x", Y288);
      $display("%x", Y289);
      $display("%x", Y290);
      $display("%x", Y291);
      $display("%x", Y292);
      $display("%x", Y293);
      $display("%x", Y294);
      $display("%x", Y295);
      $display("%x", Y296);
      $display("%x", Y297);
      $display("%x", Y298);
      $display("%x", Y299);
      $display("%x", Y300);
      $display("%x", Y301);
      $display("%x", Y302);
      $display("%x", Y303);
      $display("%x", Y304);
      $display("%x", Y305);
      $display("%x", Y306);
      $display("%x", Y307);
      $display("%x", Y308);
      $display("%x", Y309);
      $display("%x", Y310);
      $display("%x", Y311);
      $display("%x", Y312);
      $display("%x", Y313);
      $display("%x", Y314);
      $display("%x", Y315);
      $display("%x", Y316);
      $display("%x", Y317);
      $display("%x", Y318);
      $display("%x", Y319);
      $display("%x", Y320);
      $display("%x", Y321);
      $display("%x", Y322);
      $display("%x", Y323);
      $display("%x", Y324);
      $display("%x", Y325);
      $display("%x", Y326);
      $display("%x", Y327);
      $display("%x", Y328);
      $display("%x", Y329);
      $display("%x", Y330);
      $display("%x", Y331);
      $display("%x", Y332);
      $display("%x", Y333);
      $display("%x", Y334);
      $display("%x", Y335);
      $display("%x", Y336);
      $display("%x", Y337);
      $display("%x", Y338);
      $display("%x", Y339);
      $display("%x", Y340);
      $display("%x", Y341);
      $display("%x", Y342);
      $display("%x", Y343);
      $display("%x", Y344);
      $display("%x", Y345);
      $display("%x", Y346);
      $display("%x", Y347);
      $display("%x", Y348);
      $display("%x", Y349);
      $display("%x", Y350);
      $display("%x", Y351);
      $display("%x", Y352);
      $display("%x", Y353);
      $display("%x", Y354);
      $display("%x", Y355);
      $display("%x", Y356);
      $display("%x", Y357);
      $display("%x", Y358);
      $display("%x", Y359);
      $display("%x", Y360);
      $display("%x", Y361);
      $display("%x", Y362);
      $display("%x", Y363);
      $display("%x", Y364);
      $display("%x", Y365);
      $display("%x", Y366);
      $display("%x", Y367);
      $display("%x", Y368);
      $display("%x", Y369);
      $display("%x", Y370);
      $display("%x", Y371);
      $display("%x", Y372);
      $display("%x", Y373);
      $display("%x", Y374);
      $display("%x", Y375);
      $display("%x", Y376);
      $display("%x", Y377);
      $display("%x", Y378);
      $display("%x", Y379);
      $display("%x", Y380);
      $display("%x", Y381);
      $display("%x", Y382);
      $display("%x", Y383);
      $display("%x", Y384);
      $display("%x", Y385);
      $display("%x", Y386);
      $display("%x", Y387);
      $display("%x", Y388);
      $display("%x", Y389);
      $display("%x", Y390);
      $display("%x", Y391);
      $display("%x", Y392);
      $display("%x", Y393);
      $display("%x", Y394);
      $display("%x", Y395);
      $display("%x", Y396);
      $display("%x", Y397);
      $display("%x", Y398);
      $display("%x", Y399);
      $display("%x", Y400);
      $display("%x", Y401);
      $display("%x", Y402);
      $display("%x", Y403);
      $display("%x", Y404);
      $display("%x", Y405);
      $display("%x", Y406);
      $display("%x", Y407);
      $display("%x", Y408);
      $display("%x", Y409);
      $display("%x", Y410);
      $display("%x", Y411);
      $display("%x", Y412);
      $display("%x", Y413);
      $display("%x", Y414);
      $display("%x", Y415);
      $display("%x", Y416);
      $display("%x", Y417);
      $display("%x", Y418);
      $display("%x", Y419);
      $display("%x", Y420);
      $display("%x", Y421);
      $display("%x", Y422);
      $display("%x", Y423);
      $display("%x", Y424);
      $display("%x", Y425);
      $display("%x", Y426);
      $display("%x", Y427);
      $display("%x", Y428);
      $display("%x", Y429);
      $display("%x", Y430);
      $display("%x", Y431);
      $display("%x", Y432);
      $display("%x", Y433);
      $display("%x", Y434);
      $display("%x", Y435);
      $display("%x", Y436);
      $display("%x", Y437);
      $display("%x", Y438);
      $display("%x", Y439);
      $display("%x", Y440);
      $display("%x", Y441);
      $display("%x", Y442);
      $display("%x", Y443);
      $display("%x", Y444);
      $display("%x", Y445);
      $display("%x", Y446);
      $display("%x", Y447);
      $display("%x", Y448);
      $display("%x", Y449);
      $display("%x", Y450);
      $display("%x", Y451);
      $display("%x", Y452);
      $display("%x", Y453);
      $display("%x", Y454);
      $display("%x", Y455);
      $display("%x", Y456);
      $display("%x", Y457);
      $display("%x", Y458);
      $display("%x", Y459);
      $display("%x", Y460);
      $display("%x", Y461);
      $display("%x", Y462);
      $display("%x", Y463);
      $display("%x", Y464);
      $display("%x", Y465);
      $display("%x", Y466);
      $display("%x", Y467);
      $display("%x", Y468);
      $display("%x", Y469);
      $display("%x", Y470);
      $display("%x", Y471);
      $display("%x", Y472);
      $display("%x", Y473);
      $display("%x", Y474);
      $display("%x", Y475);
      $display("%x", Y476);
      $display("%x", Y477);
      $display("%x", Y478);
      $display("%x", Y479);
      $display("%x", Y480);
      $display("%x", Y481);
      $display("%x", Y482);
      $display("%x", Y483);
      $display("%x", Y484);
      $display("%x", Y485);
      $display("%x", Y486);
      $display("%x", Y487);
      $display("%x", Y488);
      $display("%x", Y489);
      $display("%x", Y490);
      $display("%x", Y491);
      $display("%x", Y492);
      $display("%x", Y493);
      $display("%x", Y494);
      $display("%x", Y495);
      $display("%x", Y496);
      $display("%x", Y497);
      $display("%x", Y498);
      $display("%x", Y499);
      $display("%x", Y500);
      $display("%x", Y501);
      $display("%x", Y502);
      $display("%x", Y503);
      $display("%x", Y504);
      $display("%x", Y505);
      $display("%x", Y506);
      $display("%x", Y507);
      $display("%x", Y508);
      $display("%x", Y509);
      $display("%x", Y510);
      $display("%x", Y511);
      $display("%x", Y512);
      $display("%x", Y513);
      $display("%x", Y514);
      $display("%x", Y515);
      $display("%x", Y516);
      $display("%x", Y517);
      $display("%x", Y518);
      $display("%x", Y519);
      $display("%x", Y520);
      $display("%x", Y521);
      $display("%x", Y522);
      $display("%x", Y523);
      $display("%x", Y524);
      $display("%x", Y525);
      $display("%x", Y526);
      $display("%x", Y527);
      $display("%x", Y528);
      $display("%x", Y529);
      $display("%x", Y530);
      $display("%x", Y531);
      $display("%x", Y532);
      $display("%x", Y533);
      $display("%x", Y534);
      $display("%x", Y535);
      $display("%x", Y536);
      $display("%x", Y537);
      $display("%x", Y538);
      $display("%x", Y539);
      $display("%x", Y540);
      $display("%x", Y541);
      $display("%x", Y542);
      $display("%x", Y543);
      $display("%x", Y544);
      $display("%x", Y545);
      $display("%x", Y546);
      $display("%x", Y547);
      $display("%x", Y548);
      $display("%x", Y549);
      $display("%x", Y550);
      $display("%x", Y551);
      $display("%x", Y552);
      $display("%x", Y553);
      $display("%x", Y554);
      $display("%x", Y555);
      $display("%x", Y556);
      $display("%x", Y557);
      $display("%x", Y558);
      $display("%x", Y559);
      $display("%x", Y560);
      $display("%x", Y561);
      $display("%x", Y562);
      $display("%x", Y563);
      $display("%x", Y564);
      $display("%x", Y565);
      $display("%x", Y566);
      $display("%x", Y567);
      $display("%x", Y568);
      $display("%x", Y569);
      $display("%x", Y570);
      $display("%x", Y571);
      $display("%x", Y572);
      $display("%x", Y573);
      $display("%x", Y574);
      $display("%x", Y575);
      $display("%x", Y576);
      $display("%x", Y577);
      $display("%x", Y578);
      $display("%x", Y579);
      $display("%x", Y580);
      $display("%x", Y581);
      $display("%x", Y582);
      $display("%x", Y583);
      $display("%x", Y584);
      $display("%x", Y585);
      $display("%x", Y586);
      $display("%x", Y587);
      $display("%x", Y588);
      $display("%x", Y589);
      $display("%x", Y590);
      $display("%x", Y591);
      $display("%x", Y592);
      $display("%x", Y593);
      $display("%x", Y594);
      $display("%x", Y595);
      $display("%x", Y596);
      $display("%x", Y597);
      $display("%x", Y598);
      $display("%x", Y599);
      $display("%x", Y600);
      $display("%x", Y601);
      $display("%x", Y602);
      $display("%x", Y603);
      $display("%x", Y604);
      $display("%x", Y605);
      $display("%x", Y606);
      $display("%x", Y607);
      $display("%x", Y608);
      $display("%x", Y609);
      $display("%x", Y610);
      $display("%x", Y611);
      $display("%x", Y612);
      $display("%x", Y613);
      $display("%x", Y614);
      $display("%x", Y615);
      $display("%x", Y616);
      $display("%x", Y617);
      $display("%x", Y618);
      $display("%x", Y619);
      $display("%x", Y620);
      $display("%x", Y621);
      $display("%x", Y622);
      $display("%x", Y623);
      $display("%x", Y624);
      $display("%x", Y625);
      $display("%x", Y626);
      $display("%x", Y627);
      $display("%x", Y628);
      $display("%x", Y629);
      $display("%x", Y630);
      $display("%x", Y631);
      $display("%x", Y632);
      $display("%x", Y633);
      $display("%x", Y634);
      $display("%x", Y635);
      $display("%x", Y636);
      $display("%x", Y637);
      $display("%x", Y638);
      $display("%x", Y639);
      $display("%x", Y640);
      $display("%x", Y641);
      $display("%x", Y642);
      $display("%x", Y643);
      $display("%x", Y644);
      $display("%x", Y645);
      $display("%x", Y646);
      $display("%x", Y647);
      $display("%x", Y648);
      $display("%x", Y649);
      $display("%x", Y650);
      $display("%x", Y651);
      $display("%x", Y652);
      $display("%x", Y653);
      $display("%x", Y654);
      $display("%x", Y655);
      $display("%x", Y656);
      $display("%x", Y657);
      $display("%x", Y658);
      $display("%x", Y659);
      $display("%x", Y660);
      $display("%x", Y661);
      $display("%x", Y662);
      $display("%x", Y663);
      $display("%x", Y664);
      $display("%x", Y665);
      $display("%x", Y666);
      $display("%x", Y667);
      $display("%x", Y668);
      $display("%x", Y669);
      $display("%x", Y670);
      $display("%x", Y671);
      $display("%x", Y672);
      $display("%x", Y673);
      $display("%x", Y674);
      $display("%x", Y675);
      $display("%x", Y676);
      $display("%x", Y677);
      $display("%x", Y678);
      $display("%x", Y679);
      $display("%x", Y680);
      $display("%x", Y681);
      $display("%x", Y682);
      $display("%x", Y683);
      $display("%x", Y684);
      $display("%x", Y685);
      $display("%x", Y686);
      $display("%x", Y687);
      $display("%x", Y688);
      $display("%x", Y689);
      $display("%x", Y690);
      $display("%x", Y691);
      $display("%x", Y692);
      $display("%x", Y693);
      $display("%x", Y694);
      $display("%x", Y695);
      $display("%x", Y696);
      $display("%x", Y697);
      $display("%x", Y698);
      $display("%x", Y699);
      $display("%x", Y700);
      $display("%x", Y701);
      $display("%x", Y702);
      $display("%x", Y703);
      $display("%x", Y704);
      $display("%x", Y705);
      $display("%x", Y706);
      $display("%x", Y707);
      $display("%x", Y708);
      $display("%x", Y709);
      $display("%x", Y710);
      $display("%x", Y711);
      $display("%x", Y712);
      $display("%x", Y713);
      $display("%x", Y714);
      $display("%x", Y715);
      $display("%x", Y716);
      $display("%x", Y717);
      $display("%x", Y718);
      $display("%x", Y719);
      $display("%x", Y720);
      $display("%x", Y721);
      $display("%x", Y722);
      $display("%x", Y723);
      $display("%x", Y724);
      $display("%x", Y725);
      $display("%x", Y726);
      $display("%x", Y727);
      $display("%x", Y728);
      $display("%x", Y729);
      $display("%x", Y730);
      $display("%x", Y731);
      $display("%x", Y732);
      $display("%x", Y733);
      $display("%x", Y734);
      $display("%x", Y735);
      $display("%x", Y736);
      $display("%x", Y737);
      $display("%x", Y738);
      $display("%x", Y739);
      $display("%x", Y740);
      $display("%x", Y741);
      $display("%x", Y742);
      $display("%x", Y743);
      $display("%x", Y744);
      $display("%x", Y745);
      $display("%x", Y746);
      $display("%x", Y747);
      $display("%x", Y748);
      $display("%x", Y749);
      $display("%x", Y750);
      $display("%x", Y751);
      $display("%x", Y752);
      $display("%x", Y753);
      $display("%x", Y754);
      $display("%x", Y755);
      $display("%x", Y756);
      $display("%x", Y757);
      $display("%x", Y758);
      $display("%x", Y759);
      $display("%x", Y760);
      $display("%x", Y761);
      $display("%x", Y762);
      $display("%x", Y763);
      $display("%x", Y764);
      $display("%x", Y765);
      $display("%x", Y766);
      $display("%x", Y767);
      $display("%x", Y768);
      $display("%x", Y769);
      $display("%x", Y770);
      $display("%x", Y771);
      $display("%x", Y772);
      $display("%x", Y773);
      $display("%x", Y774);
      $display("%x", Y775);
      $display("%x", Y776);
      $display("%x", Y777);
      $display("%x", Y778);
      $display("%x", Y779);
      $display("%x", Y780);
      $display("%x", Y781);
      $display("%x", Y782);
      $display("%x", Y783);
      $display("%x", Y784);
      $display("%x", Y785);
      $display("%x", Y786);
      $display("%x", Y787);
      $display("%x", Y788);
      $display("%x", Y789);
      $display("%x", Y790);
      $display("%x", Y791);
      $display("%x", Y792);
      $display("%x", Y793);
      $display("%x", Y794);
      $display("%x", Y795);
      $display("%x", Y796);
      $display("%x", Y797);
      $display("%x", Y798);
      $display("%x", Y799);
      $display("%x", Y800);
      $display("%x", Y801);
      $display("%x", Y802);
      $display("%x", Y803);
      $display("%x", Y804);
      $display("%x", Y805);
      $display("%x", Y806);
      $display("%x", Y807);
      $display("%x", Y808);
      $display("%x", Y809);
      $display("%x", Y810);
      $display("%x", Y811);
      $display("%x", Y812);
      $display("%x", Y813);
      $display("%x", Y814);
      $display("%x", Y815);
      $display("%x", Y816);
      $display("%x", Y817);
      $display("%x", Y818);
      $display("%x", Y819);
      $display("%x", Y820);
      $display("%x", Y821);
      $display("%x", Y822);
      $display("%x", Y823);
      $display("%x", Y824);
      $display("%x", Y825);
      $display("%x", Y826);
      $display("%x", Y827);
      $display("%x", Y828);
      $display("%x", Y829);
      $display("%x", Y830);
      $display("%x", Y831);
      $display("%x", Y832);
      $display("%x", Y833);
      $display("%x", Y834);
      $display("%x", Y835);
      $display("%x", Y836);
      $display("%x", Y837);
      $display("%x", Y838);
      $display("%x", Y839);
      $display("%x", Y840);
      $display("%x", Y841);
      $display("%x", Y842);
      $display("%x", Y843);
      $display("%x", Y844);
      $display("%x", Y845);
      $display("%x", Y846);
      $display("%x", Y847);
      $display("%x", Y848);
      $display("%x", Y849);
      $display("%x", Y850);
      $display("%x", Y851);
      $display("%x", Y852);
      $display("%x", Y853);
      $display("%x", Y854);
      $display("%x", Y855);
      $display("%x", Y856);
      $display("%x", Y857);
      $display("%x", Y858);
      $display("%x", Y859);
      $display("%x", Y860);
      $display("%x", Y861);
      $display("%x", Y862);
      $display("%x", Y863);
      $display("%x", Y864);
      $display("%x", Y865);
      $display("%x", Y866);
      $display("%x", Y867);
      $display("%x", Y868);
      $display("%x", Y869);
      $display("%x", Y870);
      $display("%x", Y871);
      $display("%x", Y872);
      $display("%x", Y873);
      $display("%x", Y874);
      $display("%x", Y875);
      $display("%x", Y876);
      $display("%x", Y877);
      $display("%x", Y878);
      $display("%x", Y879);
      $display("%x", Y880);
      $display("%x", Y881);
      $display("%x", Y882);
      $display("%x", Y883);
      $display("%x", Y884);
      $display("%x", Y885);
      $display("%x", Y886);
      $display("%x", Y887);
      $display("%x", Y888);
      $display("%x", Y889);
      $display("%x", Y890);
      $display("%x", Y891);
      $display("%x", Y892);
      $display("%x", Y893);
      $display("%x", Y894);
      $display("%x", Y895);
      $display("%x", Y896);
      $display("%x", Y897);
      $display("%x", Y898);
      $display("%x", Y899);
      $display("%x", Y900);
      $display("%x", Y901);
      $display("%x", Y902);
      $display("%x", Y903);
      $display("%x", Y904);
      $display("%x", Y905);
      $display("%x", Y906);
      $display("%x", Y907);
      $display("%x", Y908);
      $display("%x", Y909);
      $display("%x", Y910);
      $display("%x", Y911);
      $display("%x", Y912);
      $display("%x", Y913);
      $display("%x", Y914);
      $display("%x", Y915);
      $display("%x", Y916);
      $display("%x", Y917);
      $display("%x", Y918);
      $display("%x", Y919);
      $display("%x", Y920);
      $display("%x", Y921);
      $display("%x", Y922);
      $display("%x", Y923);
      $display("%x", Y924);
      $display("%x", Y925);
      $display("%x", Y926);
      $display("%x", Y927);
      $display("%x", Y928);
      $display("%x", Y929);
      $display("%x", Y930);
      $display("%x", Y931);
      $display("%x", Y932);
      $display("%x", Y933);
      $display("%x", Y934);
      $display("%x", Y935);
      $display("%x", Y936);
      $display("%x", Y937);
      $display("%x", Y938);
      $display("%x", Y939);
      $display("%x", Y940);
      $display("%x", Y941);
      $display("%x", Y942);
      $display("%x", Y943);
      $display("%x", Y944);
      $display("%x", Y945);
      $display("%x", Y946);
      $display("%x", Y947);
      $display("%x", Y948);
      $display("%x", Y949);
      $display("%x", Y950);
      $display("%x", Y951);
      $display("%x", Y952);
      $display("%x", Y953);
      $display("%x", Y954);
      $display("%x", Y955);
      $display("%x", Y956);
      $display("%x", Y957);
      $display("%x", Y958);
      $display("%x", Y959);
      $display("%x", Y960);
      $display("%x", Y961);
      $display("%x", Y962);
      $display("%x", Y963);
      $display("%x", Y964);
      $display("%x", Y965);
      $display("%x", Y966);
      $display("%x", Y967);
      $display("%x", Y968);
      $display("%x", Y969);
      $display("%x", Y970);
      $display("%x", Y971);
      $display("%x", Y972);
      $display("%x", Y973);
      $display("%x", Y974);
      $display("%x", Y975);
      $display("%x", Y976);
      $display("%x", Y977);
      $display("%x", Y978);
      $display("%x", Y979);
      $display("%x", Y980);
      $display("%x", Y981);
      $display("%x", Y982);
      $display("%x", Y983);
      $display("%x", Y984);
      $display("%x", Y985);
      $display("%x", Y986);
      $display("%x", Y987);
      $display("%x", Y988);
      $display("%x", Y989);
      $display("%x", Y990);
      $display("%x", Y991);
      $display("%x", Y992);
      $display("%x", Y993);
      $display("%x", Y994);
      $display("%x", Y995);
      $display("%x", Y996);
      $display("%x", Y997);
      $display("%x", Y998);
      $display("%x", Y999);
      $display("%x", Y1000);
      $display("%x", Y1001);
      $display("%x", Y1002);
      $display("%x", Y1003);
      $display("%x", Y1004);
      $display("%x", Y1005);
      $display("%x", Y1006);
      $display("%x", Y1007);
      $display("%x", Y1008);
      $display("%x", Y1009);
      $display("%x", Y1010);
      $display("%x", Y1011);
      $display("%x", Y1012);
      $display("%x", Y1013);
      $display("%x", Y1014);
      $display("%x", Y1015);
      $display("%x", Y1016);
      $display("%x", Y1017);
      $display("%x", Y1018);
      $display("%x", Y1019);
      $display("%x", Y1020);
      $display("%x", Y1021);
      $display("%x", Y1022);
      $display("%x", Y1023);
      // Wait until next_out goes high, then wait one clock cycle and begin receiving data
      @(posedge next_out);
      @(posedge clk); #1;
      $display("--- begin output 2---");

      for (m=0; m < 0; m=m+1) begin
         $display("%x", Y0);
         $display("%x", Y1);
         $display("%x", Y2);
         $display("%x", Y3);
         $display("%x", Y4);
         $display("%x", Y5);
         $display("%x", Y6);
         $display("%x", Y7);
         $display("%x", Y8);
         $display("%x", Y9);
         $display("%x", Y10);
         $display("%x", Y11);
         $display("%x", Y12);
         $display("%x", Y13);
         $display("%x", Y14);
         $display("%x", Y15);
         $display("%x", Y16);
         $display("%x", Y17);
         $display("%x", Y18);
         $display("%x", Y19);
         $display("%x", Y20);
         $display("%x", Y21);
         $display("%x", Y22);
         $display("%x", Y23);
         $display("%x", Y24);
         $display("%x", Y25);
         $display("%x", Y26);
         $display("%x", Y27);
         $display("%x", Y28);
         $display("%x", Y29);
         $display("%x", Y30);
         $display("%x", Y31);
         $display("%x", Y32);
         $display("%x", Y33);
         $display("%x", Y34);
         $display("%x", Y35);
         $display("%x", Y36);
         $display("%x", Y37);
         $display("%x", Y38);
         $display("%x", Y39);
         $display("%x", Y40);
         $display("%x", Y41);
         $display("%x", Y42);
         $display("%x", Y43);
         $display("%x", Y44);
         $display("%x", Y45);
         $display("%x", Y46);
         $display("%x", Y47);
         $display("%x", Y48);
         $display("%x", Y49);
         $display("%x", Y50);
         $display("%x", Y51);
         $display("%x", Y52);
         $display("%x", Y53);
         $display("%x", Y54);
         $display("%x", Y55);
         $display("%x", Y56);
         $display("%x", Y57);
         $display("%x", Y58);
         $display("%x", Y59);
         $display("%x", Y60);
         $display("%x", Y61);
         $display("%x", Y62);
         $display("%x", Y63);
         $display("%x", Y64);
         $display("%x", Y65);
         $display("%x", Y66);
         $display("%x", Y67);
         $display("%x", Y68);
         $display("%x", Y69);
         $display("%x", Y70);
         $display("%x", Y71);
         $display("%x", Y72);
         $display("%x", Y73);
         $display("%x", Y74);
         $display("%x", Y75);
         $display("%x", Y76);
         $display("%x", Y77);
         $display("%x", Y78);
         $display("%x", Y79);
         $display("%x", Y80);
         $display("%x", Y81);
         $display("%x", Y82);
         $display("%x", Y83);
         $display("%x", Y84);
         $display("%x", Y85);
         $display("%x", Y86);
         $display("%x", Y87);
         $display("%x", Y88);
         $display("%x", Y89);
         $display("%x", Y90);
         $display("%x", Y91);
         $display("%x", Y92);
         $display("%x", Y93);
         $display("%x", Y94);
         $display("%x", Y95);
         $display("%x", Y96);
         $display("%x", Y97);
         $display("%x", Y98);
         $display("%x", Y99);
         $display("%x", Y100);
         $display("%x", Y101);
         $display("%x", Y102);
         $display("%x", Y103);
         $display("%x", Y104);
         $display("%x", Y105);
         $display("%x", Y106);
         $display("%x", Y107);
         $display("%x", Y108);
         $display("%x", Y109);
         $display("%x", Y110);
         $display("%x", Y111);
         $display("%x", Y112);
         $display("%x", Y113);
         $display("%x", Y114);
         $display("%x", Y115);
         $display("%x", Y116);
         $display("%x", Y117);
         $display("%x", Y118);
         $display("%x", Y119);
         $display("%x", Y120);
         $display("%x", Y121);
         $display("%x", Y122);
         $display("%x", Y123);
         $display("%x", Y124);
         $display("%x", Y125);
         $display("%x", Y126);
         $display("%x", Y127);
         $display("%x", Y128);
         $display("%x", Y129);
         $display("%x", Y130);
         $display("%x", Y131);
         $display("%x", Y132);
         $display("%x", Y133);
         $display("%x", Y134);
         $display("%x", Y135);
         $display("%x", Y136);
         $display("%x", Y137);
         $display("%x", Y138);
         $display("%x", Y139);
         $display("%x", Y140);
         $display("%x", Y141);
         $display("%x", Y142);
         $display("%x", Y143);
         $display("%x", Y144);
         $display("%x", Y145);
         $display("%x", Y146);
         $display("%x", Y147);
         $display("%x", Y148);
         $display("%x", Y149);
         $display("%x", Y150);
         $display("%x", Y151);
         $display("%x", Y152);
         $display("%x", Y153);
         $display("%x", Y154);
         $display("%x", Y155);
         $display("%x", Y156);
         $display("%x", Y157);
         $display("%x", Y158);
         $display("%x", Y159);
         $display("%x", Y160);
         $display("%x", Y161);
         $display("%x", Y162);
         $display("%x", Y163);
         $display("%x", Y164);
         $display("%x", Y165);
         $display("%x", Y166);
         $display("%x", Y167);
         $display("%x", Y168);
         $display("%x", Y169);
         $display("%x", Y170);
         $display("%x", Y171);
         $display("%x", Y172);
         $display("%x", Y173);
         $display("%x", Y174);
         $display("%x", Y175);
         $display("%x", Y176);
         $display("%x", Y177);
         $display("%x", Y178);
         $display("%x", Y179);
         $display("%x", Y180);
         $display("%x", Y181);
         $display("%x", Y182);
         $display("%x", Y183);
         $display("%x", Y184);
         $display("%x", Y185);
         $display("%x", Y186);
         $display("%x", Y187);
         $display("%x", Y188);
         $display("%x", Y189);
         $display("%x", Y190);
         $display("%x", Y191);
         $display("%x", Y192);
         $display("%x", Y193);
         $display("%x", Y194);
         $display("%x", Y195);
         $display("%x", Y196);
         $display("%x", Y197);
         $display("%x", Y198);
         $display("%x", Y199);
         $display("%x", Y200);
         $display("%x", Y201);
         $display("%x", Y202);
         $display("%x", Y203);
         $display("%x", Y204);
         $display("%x", Y205);
         $display("%x", Y206);
         $display("%x", Y207);
         $display("%x", Y208);
         $display("%x", Y209);
         $display("%x", Y210);
         $display("%x", Y211);
         $display("%x", Y212);
         $display("%x", Y213);
         $display("%x", Y214);
         $display("%x", Y215);
         $display("%x", Y216);
         $display("%x", Y217);
         $display("%x", Y218);
         $display("%x", Y219);
         $display("%x", Y220);
         $display("%x", Y221);
         $display("%x", Y222);
         $display("%x", Y223);
         $display("%x", Y224);
         $display("%x", Y225);
         $display("%x", Y226);
         $display("%x", Y227);
         $display("%x", Y228);
         $display("%x", Y229);
         $display("%x", Y230);
         $display("%x", Y231);
         $display("%x", Y232);
         $display("%x", Y233);
         $display("%x", Y234);
         $display("%x", Y235);
         $display("%x", Y236);
         $display("%x", Y237);
         $display("%x", Y238);
         $display("%x", Y239);
         $display("%x", Y240);
         $display("%x", Y241);
         $display("%x", Y242);
         $display("%x", Y243);
         $display("%x", Y244);
         $display("%x", Y245);
         $display("%x", Y246);
         $display("%x", Y247);
         $display("%x", Y248);
         $display("%x", Y249);
         $display("%x", Y250);
         $display("%x", Y251);
         $display("%x", Y252);
         $display("%x", Y253);
         $display("%x", Y254);
         $display("%x", Y255);
         $display("%x", Y256);
         $display("%x", Y257);
         $display("%x", Y258);
         $display("%x", Y259);
         $display("%x", Y260);
         $display("%x", Y261);
         $display("%x", Y262);
         $display("%x", Y263);
         $display("%x", Y264);
         $display("%x", Y265);
         $display("%x", Y266);
         $display("%x", Y267);
         $display("%x", Y268);
         $display("%x", Y269);
         $display("%x", Y270);
         $display("%x", Y271);
         $display("%x", Y272);
         $display("%x", Y273);
         $display("%x", Y274);
         $display("%x", Y275);
         $display("%x", Y276);
         $display("%x", Y277);
         $display("%x", Y278);
         $display("%x", Y279);
         $display("%x", Y280);
         $display("%x", Y281);
         $display("%x", Y282);
         $display("%x", Y283);
         $display("%x", Y284);
         $display("%x", Y285);
         $display("%x", Y286);
         $display("%x", Y287);
         $display("%x", Y288);
         $display("%x", Y289);
         $display("%x", Y290);
         $display("%x", Y291);
         $display("%x", Y292);
         $display("%x", Y293);
         $display("%x", Y294);
         $display("%x", Y295);
         $display("%x", Y296);
         $display("%x", Y297);
         $display("%x", Y298);
         $display("%x", Y299);
         $display("%x", Y300);
         $display("%x", Y301);
         $display("%x", Y302);
         $display("%x", Y303);
         $display("%x", Y304);
         $display("%x", Y305);
         $display("%x", Y306);
         $display("%x", Y307);
         $display("%x", Y308);
         $display("%x", Y309);
         $display("%x", Y310);
         $display("%x", Y311);
         $display("%x", Y312);
         $display("%x", Y313);
         $display("%x", Y314);
         $display("%x", Y315);
         $display("%x", Y316);
         $display("%x", Y317);
         $display("%x", Y318);
         $display("%x", Y319);
         $display("%x", Y320);
         $display("%x", Y321);
         $display("%x", Y322);
         $display("%x", Y323);
         $display("%x", Y324);
         $display("%x", Y325);
         $display("%x", Y326);
         $display("%x", Y327);
         $display("%x", Y328);
         $display("%x", Y329);
         $display("%x", Y330);
         $display("%x", Y331);
         $display("%x", Y332);
         $display("%x", Y333);
         $display("%x", Y334);
         $display("%x", Y335);
         $display("%x", Y336);
         $display("%x", Y337);
         $display("%x", Y338);
         $display("%x", Y339);
         $display("%x", Y340);
         $display("%x", Y341);
         $display("%x", Y342);
         $display("%x", Y343);
         $display("%x", Y344);
         $display("%x", Y345);
         $display("%x", Y346);
         $display("%x", Y347);
         $display("%x", Y348);
         $display("%x", Y349);
         $display("%x", Y350);
         $display("%x", Y351);
         $display("%x", Y352);
         $display("%x", Y353);
         $display("%x", Y354);
         $display("%x", Y355);
         $display("%x", Y356);
         $display("%x", Y357);
         $display("%x", Y358);
         $display("%x", Y359);
         $display("%x", Y360);
         $display("%x", Y361);
         $display("%x", Y362);
         $display("%x", Y363);
         $display("%x", Y364);
         $display("%x", Y365);
         $display("%x", Y366);
         $display("%x", Y367);
         $display("%x", Y368);
         $display("%x", Y369);
         $display("%x", Y370);
         $display("%x", Y371);
         $display("%x", Y372);
         $display("%x", Y373);
         $display("%x", Y374);
         $display("%x", Y375);
         $display("%x", Y376);
         $display("%x", Y377);
         $display("%x", Y378);
         $display("%x", Y379);
         $display("%x", Y380);
         $display("%x", Y381);
         $display("%x", Y382);
         $display("%x", Y383);
         $display("%x", Y384);
         $display("%x", Y385);
         $display("%x", Y386);
         $display("%x", Y387);
         $display("%x", Y388);
         $display("%x", Y389);
         $display("%x", Y390);
         $display("%x", Y391);
         $display("%x", Y392);
         $display("%x", Y393);
         $display("%x", Y394);
         $display("%x", Y395);
         $display("%x", Y396);
         $display("%x", Y397);
         $display("%x", Y398);
         $display("%x", Y399);
         $display("%x", Y400);
         $display("%x", Y401);
         $display("%x", Y402);
         $display("%x", Y403);
         $display("%x", Y404);
         $display("%x", Y405);
         $display("%x", Y406);
         $display("%x", Y407);
         $display("%x", Y408);
         $display("%x", Y409);
         $display("%x", Y410);
         $display("%x", Y411);
         $display("%x", Y412);
         $display("%x", Y413);
         $display("%x", Y414);
         $display("%x", Y415);
         $display("%x", Y416);
         $display("%x", Y417);
         $display("%x", Y418);
         $display("%x", Y419);
         $display("%x", Y420);
         $display("%x", Y421);
         $display("%x", Y422);
         $display("%x", Y423);
         $display("%x", Y424);
         $display("%x", Y425);
         $display("%x", Y426);
         $display("%x", Y427);
         $display("%x", Y428);
         $display("%x", Y429);
         $display("%x", Y430);
         $display("%x", Y431);
         $display("%x", Y432);
         $display("%x", Y433);
         $display("%x", Y434);
         $display("%x", Y435);
         $display("%x", Y436);
         $display("%x", Y437);
         $display("%x", Y438);
         $display("%x", Y439);
         $display("%x", Y440);
         $display("%x", Y441);
         $display("%x", Y442);
         $display("%x", Y443);
         $display("%x", Y444);
         $display("%x", Y445);
         $display("%x", Y446);
         $display("%x", Y447);
         $display("%x", Y448);
         $display("%x", Y449);
         $display("%x", Y450);
         $display("%x", Y451);
         $display("%x", Y452);
         $display("%x", Y453);
         $display("%x", Y454);
         $display("%x", Y455);
         $display("%x", Y456);
         $display("%x", Y457);
         $display("%x", Y458);
         $display("%x", Y459);
         $display("%x", Y460);
         $display("%x", Y461);
         $display("%x", Y462);
         $display("%x", Y463);
         $display("%x", Y464);
         $display("%x", Y465);
         $display("%x", Y466);
         $display("%x", Y467);
         $display("%x", Y468);
         $display("%x", Y469);
         $display("%x", Y470);
         $display("%x", Y471);
         $display("%x", Y472);
         $display("%x", Y473);
         $display("%x", Y474);
         $display("%x", Y475);
         $display("%x", Y476);
         $display("%x", Y477);
         $display("%x", Y478);
         $display("%x", Y479);
         $display("%x", Y480);
         $display("%x", Y481);
         $display("%x", Y482);
         $display("%x", Y483);
         $display("%x", Y484);
         $display("%x", Y485);
         $display("%x", Y486);
         $display("%x", Y487);
         $display("%x", Y488);
         $display("%x", Y489);
         $display("%x", Y490);
         $display("%x", Y491);
         $display("%x", Y492);
         $display("%x", Y493);
         $display("%x", Y494);
         $display("%x", Y495);
         $display("%x", Y496);
         $display("%x", Y497);
         $display("%x", Y498);
         $display("%x", Y499);
         $display("%x", Y500);
         $display("%x", Y501);
         $display("%x", Y502);
         $display("%x", Y503);
         $display("%x", Y504);
         $display("%x", Y505);
         $display("%x", Y506);
         $display("%x", Y507);
         $display("%x", Y508);
         $display("%x", Y509);
         $display("%x", Y510);
         $display("%x", Y511);
         $display("%x", Y512);
         $display("%x", Y513);
         $display("%x", Y514);
         $display("%x", Y515);
         $display("%x", Y516);
         $display("%x", Y517);
         $display("%x", Y518);
         $display("%x", Y519);
         $display("%x", Y520);
         $display("%x", Y521);
         $display("%x", Y522);
         $display("%x", Y523);
         $display("%x", Y524);
         $display("%x", Y525);
         $display("%x", Y526);
         $display("%x", Y527);
         $display("%x", Y528);
         $display("%x", Y529);
         $display("%x", Y530);
         $display("%x", Y531);
         $display("%x", Y532);
         $display("%x", Y533);
         $display("%x", Y534);
         $display("%x", Y535);
         $display("%x", Y536);
         $display("%x", Y537);
         $display("%x", Y538);
         $display("%x", Y539);
         $display("%x", Y540);
         $display("%x", Y541);
         $display("%x", Y542);
         $display("%x", Y543);
         $display("%x", Y544);
         $display("%x", Y545);
         $display("%x", Y546);
         $display("%x", Y547);
         $display("%x", Y548);
         $display("%x", Y549);
         $display("%x", Y550);
         $display("%x", Y551);
         $display("%x", Y552);
         $display("%x", Y553);
         $display("%x", Y554);
         $display("%x", Y555);
         $display("%x", Y556);
         $display("%x", Y557);
         $display("%x", Y558);
         $display("%x", Y559);
         $display("%x", Y560);
         $display("%x", Y561);
         $display("%x", Y562);
         $display("%x", Y563);
         $display("%x", Y564);
         $display("%x", Y565);
         $display("%x", Y566);
         $display("%x", Y567);
         $display("%x", Y568);
         $display("%x", Y569);
         $display("%x", Y570);
         $display("%x", Y571);
         $display("%x", Y572);
         $display("%x", Y573);
         $display("%x", Y574);
         $display("%x", Y575);
         $display("%x", Y576);
         $display("%x", Y577);
         $display("%x", Y578);
         $display("%x", Y579);
         $display("%x", Y580);
         $display("%x", Y581);
         $display("%x", Y582);
         $display("%x", Y583);
         $display("%x", Y584);
         $display("%x", Y585);
         $display("%x", Y586);
         $display("%x", Y587);
         $display("%x", Y588);
         $display("%x", Y589);
         $display("%x", Y590);
         $display("%x", Y591);
         $display("%x", Y592);
         $display("%x", Y593);
         $display("%x", Y594);
         $display("%x", Y595);
         $display("%x", Y596);
         $display("%x", Y597);
         $display("%x", Y598);
         $display("%x", Y599);
         $display("%x", Y600);
         $display("%x", Y601);
         $display("%x", Y602);
         $display("%x", Y603);
         $display("%x", Y604);
         $display("%x", Y605);
         $display("%x", Y606);
         $display("%x", Y607);
         $display("%x", Y608);
         $display("%x", Y609);
         $display("%x", Y610);
         $display("%x", Y611);
         $display("%x", Y612);
         $display("%x", Y613);
         $display("%x", Y614);
         $display("%x", Y615);
         $display("%x", Y616);
         $display("%x", Y617);
         $display("%x", Y618);
         $display("%x", Y619);
         $display("%x", Y620);
         $display("%x", Y621);
         $display("%x", Y622);
         $display("%x", Y623);
         $display("%x", Y624);
         $display("%x", Y625);
         $display("%x", Y626);
         $display("%x", Y627);
         $display("%x", Y628);
         $display("%x", Y629);
         $display("%x", Y630);
         $display("%x", Y631);
         $display("%x", Y632);
         $display("%x", Y633);
         $display("%x", Y634);
         $display("%x", Y635);
         $display("%x", Y636);
         $display("%x", Y637);
         $display("%x", Y638);
         $display("%x", Y639);
         $display("%x", Y640);
         $display("%x", Y641);
         $display("%x", Y642);
         $display("%x", Y643);
         $display("%x", Y644);
         $display("%x", Y645);
         $display("%x", Y646);
         $display("%x", Y647);
         $display("%x", Y648);
         $display("%x", Y649);
         $display("%x", Y650);
         $display("%x", Y651);
         $display("%x", Y652);
         $display("%x", Y653);
         $display("%x", Y654);
         $display("%x", Y655);
         $display("%x", Y656);
         $display("%x", Y657);
         $display("%x", Y658);
         $display("%x", Y659);
         $display("%x", Y660);
         $display("%x", Y661);
         $display("%x", Y662);
         $display("%x", Y663);
         $display("%x", Y664);
         $display("%x", Y665);
         $display("%x", Y666);
         $display("%x", Y667);
         $display("%x", Y668);
         $display("%x", Y669);
         $display("%x", Y670);
         $display("%x", Y671);
         $display("%x", Y672);
         $display("%x", Y673);
         $display("%x", Y674);
         $display("%x", Y675);
         $display("%x", Y676);
         $display("%x", Y677);
         $display("%x", Y678);
         $display("%x", Y679);
         $display("%x", Y680);
         $display("%x", Y681);
         $display("%x", Y682);
         $display("%x", Y683);
         $display("%x", Y684);
         $display("%x", Y685);
         $display("%x", Y686);
         $display("%x", Y687);
         $display("%x", Y688);
         $display("%x", Y689);
         $display("%x", Y690);
         $display("%x", Y691);
         $display("%x", Y692);
         $display("%x", Y693);
         $display("%x", Y694);
         $display("%x", Y695);
         $display("%x", Y696);
         $display("%x", Y697);
         $display("%x", Y698);
         $display("%x", Y699);
         $display("%x", Y700);
         $display("%x", Y701);
         $display("%x", Y702);
         $display("%x", Y703);
         $display("%x", Y704);
         $display("%x", Y705);
         $display("%x", Y706);
         $display("%x", Y707);
         $display("%x", Y708);
         $display("%x", Y709);
         $display("%x", Y710);
         $display("%x", Y711);
         $display("%x", Y712);
         $display("%x", Y713);
         $display("%x", Y714);
         $display("%x", Y715);
         $display("%x", Y716);
         $display("%x", Y717);
         $display("%x", Y718);
         $display("%x", Y719);
         $display("%x", Y720);
         $display("%x", Y721);
         $display("%x", Y722);
         $display("%x", Y723);
         $display("%x", Y724);
         $display("%x", Y725);
         $display("%x", Y726);
         $display("%x", Y727);
         $display("%x", Y728);
         $display("%x", Y729);
         $display("%x", Y730);
         $display("%x", Y731);
         $display("%x", Y732);
         $display("%x", Y733);
         $display("%x", Y734);
         $display("%x", Y735);
         $display("%x", Y736);
         $display("%x", Y737);
         $display("%x", Y738);
         $display("%x", Y739);
         $display("%x", Y740);
         $display("%x", Y741);
         $display("%x", Y742);
         $display("%x", Y743);
         $display("%x", Y744);
         $display("%x", Y745);
         $display("%x", Y746);
         $display("%x", Y747);
         $display("%x", Y748);
         $display("%x", Y749);
         $display("%x", Y750);
         $display("%x", Y751);
         $display("%x", Y752);
         $display("%x", Y753);
         $display("%x", Y754);
         $display("%x", Y755);
         $display("%x", Y756);
         $display("%x", Y757);
         $display("%x", Y758);
         $display("%x", Y759);
         $display("%x", Y760);
         $display("%x", Y761);
         $display("%x", Y762);
         $display("%x", Y763);
         $display("%x", Y764);
         $display("%x", Y765);
         $display("%x", Y766);
         $display("%x", Y767);
         $display("%x", Y768);
         $display("%x", Y769);
         $display("%x", Y770);
         $display("%x", Y771);
         $display("%x", Y772);
         $display("%x", Y773);
         $display("%x", Y774);
         $display("%x", Y775);
         $display("%x", Y776);
         $display("%x", Y777);
         $display("%x", Y778);
         $display("%x", Y779);
         $display("%x", Y780);
         $display("%x", Y781);
         $display("%x", Y782);
         $display("%x", Y783);
         $display("%x", Y784);
         $display("%x", Y785);
         $display("%x", Y786);
         $display("%x", Y787);
         $display("%x", Y788);
         $display("%x", Y789);
         $display("%x", Y790);
         $display("%x", Y791);
         $display("%x", Y792);
         $display("%x", Y793);
         $display("%x", Y794);
         $display("%x", Y795);
         $display("%x", Y796);
         $display("%x", Y797);
         $display("%x", Y798);
         $display("%x", Y799);
         $display("%x", Y800);
         $display("%x", Y801);
         $display("%x", Y802);
         $display("%x", Y803);
         $display("%x", Y804);
         $display("%x", Y805);
         $display("%x", Y806);
         $display("%x", Y807);
         $display("%x", Y808);
         $display("%x", Y809);
         $display("%x", Y810);
         $display("%x", Y811);
         $display("%x", Y812);
         $display("%x", Y813);
         $display("%x", Y814);
         $display("%x", Y815);
         $display("%x", Y816);
         $display("%x", Y817);
         $display("%x", Y818);
         $display("%x", Y819);
         $display("%x", Y820);
         $display("%x", Y821);
         $display("%x", Y822);
         $display("%x", Y823);
         $display("%x", Y824);
         $display("%x", Y825);
         $display("%x", Y826);
         $display("%x", Y827);
         $display("%x", Y828);
         $display("%x", Y829);
         $display("%x", Y830);
         $display("%x", Y831);
         $display("%x", Y832);
         $display("%x", Y833);
         $display("%x", Y834);
         $display("%x", Y835);
         $display("%x", Y836);
         $display("%x", Y837);
         $display("%x", Y838);
         $display("%x", Y839);
         $display("%x", Y840);
         $display("%x", Y841);
         $display("%x", Y842);
         $display("%x", Y843);
         $display("%x", Y844);
         $display("%x", Y845);
         $display("%x", Y846);
         $display("%x", Y847);
         $display("%x", Y848);
         $display("%x", Y849);
         $display("%x", Y850);
         $display("%x", Y851);
         $display("%x", Y852);
         $display("%x", Y853);
         $display("%x", Y854);
         $display("%x", Y855);
         $display("%x", Y856);
         $display("%x", Y857);
         $display("%x", Y858);
         $display("%x", Y859);
         $display("%x", Y860);
         $display("%x", Y861);
         $display("%x", Y862);
         $display("%x", Y863);
         $display("%x", Y864);
         $display("%x", Y865);
         $display("%x", Y866);
         $display("%x", Y867);
         $display("%x", Y868);
         $display("%x", Y869);
         $display("%x", Y870);
         $display("%x", Y871);
         $display("%x", Y872);
         $display("%x", Y873);
         $display("%x", Y874);
         $display("%x", Y875);
         $display("%x", Y876);
         $display("%x", Y877);
         $display("%x", Y878);
         $display("%x", Y879);
         $display("%x", Y880);
         $display("%x", Y881);
         $display("%x", Y882);
         $display("%x", Y883);
         $display("%x", Y884);
         $display("%x", Y885);
         $display("%x", Y886);
         $display("%x", Y887);
         $display("%x", Y888);
         $display("%x", Y889);
         $display("%x", Y890);
         $display("%x", Y891);
         $display("%x", Y892);
         $display("%x", Y893);
         $display("%x", Y894);
         $display("%x", Y895);
         $display("%x", Y896);
         $display("%x", Y897);
         $display("%x", Y898);
         $display("%x", Y899);
         $display("%x", Y900);
         $display("%x", Y901);
         $display("%x", Y902);
         $display("%x", Y903);
         $display("%x", Y904);
         $display("%x", Y905);
         $display("%x", Y906);
         $display("%x", Y907);
         $display("%x", Y908);
         $display("%x", Y909);
         $display("%x", Y910);
         $display("%x", Y911);
         $display("%x", Y912);
         $display("%x", Y913);
         $display("%x", Y914);
         $display("%x", Y915);
         $display("%x", Y916);
         $display("%x", Y917);
         $display("%x", Y918);
         $display("%x", Y919);
         $display("%x", Y920);
         $display("%x", Y921);
         $display("%x", Y922);
         $display("%x", Y923);
         $display("%x", Y924);
         $display("%x", Y925);
         $display("%x", Y926);
         $display("%x", Y927);
         $display("%x", Y928);
         $display("%x", Y929);
         $display("%x", Y930);
         $display("%x", Y931);
         $display("%x", Y932);
         $display("%x", Y933);
         $display("%x", Y934);
         $display("%x", Y935);
         $display("%x", Y936);
         $display("%x", Y937);
         $display("%x", Y938);
         $display("%x", Y939);
         $display("%x", Y940);
         $display("%x", Y941);
         $display("%x", Y942);
         $display("%x", Y943);
         $display("%x", Y944);
         $display("%x", Y945);
         $display("%x", Y946);
         $display("%x", Y947);
         $display("%x", Y948);
         $display("%x", Y949);
         $display("%x", Y950);
         $display("%x", Y951);
         $display("%x", Y952);
         $display("%x", Y953);
         $display("%x", Y954);
         $display("%x", Y955);
         $display("%x", Y956);
         $display("%x", Y957);
         $display("%x", Y958);
         $display("%x", Y959);
         $display("%x", Y960);
         $display("%x", Y961);
         $display("%x", Y962);
         $display("%x", Y963);
         $display("%x", Y964);
         $display("%x", Y965);
         $display("%x", Y966);
         $display("%x", Y967);
         $display("%x", Y968);
         $display("%x", Y969);
         $display("%x", Y970);
         $display("%x", Y971);
         $display("%x", Y972);
         $display("%x", Y973);
         $display("%x", Y974);
         $display("%x", Y975);
         $display("%x", Y976);
         $display("%x", Y977);
         $display("%x", Y978);
         $display("%x", Y979);
         $display("%x", Y980);
         $display("%x", Y981);
         $display("%x", Y982);
         $display("%x", Y983);
         $display("%x", Y984);
         $display("%x", Y985);
         $display("%x", Y986);
         $display("%x", Y987);
         $display("%x", Y988);
         $display("%x", Y989);
         $display("%x", Y990);
         $display("%x", Y991);
         $display("%x", Y992);
         $display("%x", Y993);
         $display("%x", Y994);
         $display("%x", Y995);
         $display("%x", Y996);
         $display("%x", Y997);
         $display("%x", Y998);
         $display("%x", Y999);
         $display("%x", Y1000);
         $display("%x", Y1001);
         $display("%x", Y1002);
         $display("%x", Y1003);
         $display("%x", Y1004);
         $display("%x", Y1005);
         $display("%x", Y1006);
         $display("%x", Y1007);
         $display("%x", Y1008);
         $display("%x", Y1009);
         $display("%x", Y1010);
         $display("%x", Y1011);
         $display("%x", Y1012);
         $display("%x", Y1013);
         $display("%x", Y1014);
         $display("%x", Y1015);
         $display("%x", Y1016);
         $display("%x", Y1017);
         $display("%x", Y1018);
         $display("%x", Y1019);
         $display("%x", Y1020);
         $display("%x", Y1021);
         $display("%x", Y1022);
         $display("%x", Y1023);
         @(posedge clk); #1;
      end
      $display("%x", Y0);
      $display("%x", Y1);
      $display("%x", Y2);
      $display("%x", Y3);
      $display("%x", Y4);
      $display("%x", Y5);
      $display("%x", Y6);
      $display("%x", Y7);
      $display("%x", Y8);
      $display("%x", Y9);
      $display("%x", Y10);
      $display("%x", Y11);
      $display("%x", Y12);
      $display("%x", Y13);
      $display("%x", Y14);
      $display("%x", Y15);
      $display("%x", Y16);
      $display("%x", Y17);
      $display("%x", Y18);
      $display("%x", Y19);
      $display("%x", Y20);
      $display("%x", Y21);
      $display("%x", Y22);
      $display("%x", Y23);
      $display("%x", Y24);
      $display("%x", Y25);
      $display("%x", Y26);
      $display("%x", Y27);
      $display("%x", Y28);
      $display("%x", Y29);
      $display("%x", Y30);
      $display("%x", Y31);
      $display("%x", Y32);
      $display("%x", Y33);
      $display("%x", Y34);
      $display("%x", Y35);
      $display("%x", Y36);
      $display("%x", Y37);
      $display("%x", Y38);
      $display("%x", Y39);
      $display("%x", Y40);
      $display("%x", Y41);
      $display("%x", Y42);
      $display("%x", Y43);
      $display("%x", Y44);
      $display("%x", Y45);
      $display("%x", Y46);
      $display("%x", Y47);
      $display("%x", Y48);
      $display("%x", Y49);
      $display("%x", Y50);
      $display("%x", Y51);
      $display("%x", Y52);
      $display("%x", Y53);
      $display("%x", Y54);
      $display("%x", Y55);
      $display("%x", Y56);
      $display("%x", Y57);
      $display("%x", Y58);
      $display("%x", Y59);
      $display("%x", Y60);
      $display("%x", Y61);
      $display("%x", Y62);
      $display("%x", Y63);
      $display("%x", Y64);
      $display("%x", Y65);
      $display("%x", Y66);
      $display("%x", Y67);
      $display("%x", Y68);
      $display("%x", Y69);
      $display("%x", Y70);
      $display("%x", Y71);
      $display("%x", Y72);
      $display("%x", Y73);
      $display("%x", Y74);
      $display("%x", Y75);
      $display("%x", Y76);
      $display("%x", Y77);
      $display("%x", Y78);
      $display("%x", Y79);
      $display("%x", Y80);
      $display("%x", Y81);
      $display("%x", Y82);
      $display("%x", Y83);
      $display("%x", Y84);
      $display("%x", Y85);
      $display("%x", Y86);
      $display("%x", Y87);
      $display("%x", Y88);
      $display("%x", Y89);
      $display("%x", Y90);
      $display("%x", Y91);
      $display("%x", Y92);
      $display("%x", Y93);
      $display("%x", Y94);
      $display("%x", Y95);
      $display("%x", Y96);
      $display("%x", Y97);
      $display("%x", Y98);
      $display("%x", Y99);
      $display("%x", Y100);
      $display("%x", Y101);
      $display("%x", Y102);
      $display("%x", Y103);
      $display("%x", Y104);
      $display("%x", Y105);
      $display("%x", Y106);
      $display("%x", Y107);
      $display("%x", Y108);
      $display("%x", Y109);
      $display("%x", Y110);
      $display("%x", Y111);
      $display("%x", Y112);
      $display("%x", Y113);
      $display("%x", Y114);
      $display("%x", Y115);
      $display("%x", Y116);
      $display("%x", Y117);
      $display("%x", Y118);
      $display("%x", Y119);
      $display("%x", Y120);
      $display("%x", Y121);
      $display("%x", Y122);
      $display("%x", Y123);
      $display("%x", Y124);
      $display("%x", Y125);
      $display("%x", Y126);
      $display("%x", Y127);
      $display("%x", Y128);
      $display("%x", Y129);
      $display("%x", Y130);
      $display("%x", Y131);
      $display("%x", Y132);
      $display("%x", Y133);
      $display("%x", Y134);
      $display("%x", Y135);
      $display("%x", Y136);
      $display("%x", Y137);
      $display("%x", Y138);
      $display("%x", Y139);
      $display("%x", Y140);
      $display("%x", Y141);
      $display("%x", Y142);
      $display("%x", Y143);
      $display("%x", Y144);
      $display("%x", Y145);
      $display("%x", Y146);
      $display("%x", Y147);
      $display("%x", Y148);
      $display("%x", Y149);
      $display("%x", Y150);
      $display("%x", Y151);
      $display("%x", Y152);
      $display("%x", Y153);
      $display("%x", Y154);
      $display("%x", Y155);
      $display("%x", Y156);
      $display("%x", Y157);
      $display("%x", Y158);
      $display("%x", Y159);
      $display("%x", Y160);
      $display("%x", Y161);
      $display("%x", Y162);
      $display("%x", Y163);
      $display("%x", Y164);
      $display("%x", Y165);
      $display("%x", Y166);
      $display("%x", Y167);
      $display("%x", Y168);
      $display("%x", Y169);
      $display("%x", Y170);
      $display("%x", Y171);
      $display("%x", Y172);
      $display("%x", Y173);
      $display("%x", Y174);
      $display("%x", Y175);
      $display("%x", Y176);
      $display("%x", Y177);
      $display("%x", Y178);
      $display("%x", Y179);
      $display("%x", Y180);
      $display("%x", Y181);
      $display("%x", Y182);
      $display("%x", Y183);
      $display("%x", Y184);
      $display("%x", Y185);
      $display("%x", Y186);
      $display("%x", Y187);
      $display("%x", Y188);
      $display("%x", Y189);
      $display("%x", Y190);
      $display("%x", Y191);
      $display("%x", Y192);
      $display("%x", Y193);
      $display("%x", Y194);
      $display("%x", Y195);
      $display("%x", Y196);
      $display("%x", Y197);
      $display("%x", Y198);
      $display("%x", Y199);
      $display("%x", Y200);
      $display("%x", Y201);
      $display("%x", Y202);
      $display("%x", Y203);
      $display("%x", Y204);
      $display("%x", Y205);
      $display("%x", Y206);
      $display("%x", Y207);
      $display("%x", Y208);
      $display("%x", Y209);
      $display("%x", Y210);
      $display("%x", Y211);
      $display("%x", Y212);
      $display("%x", Y213);
      $display("%x", Y214);
      $display("%x", Y215);
      $display("%x", Y216);
      $display("%x", Y217);
      $display("%x", Y218);
      $display("%x", Y219);
      $display("%x", Y220);
      $display("%x", Y221);
      $display("%x", Y222);
      $display("%x", Y223);
      $display("%x", Y224);
      $display("%x", Y225);
      $display("%x", Y226);
      $display("%x", Y227);
      $display("%x", Y228);
      $display("%x", Y229);
      $display("%x", Y230);
      $display("%x", Y231);
      $display("%x", Y232);
      $display("%x", Y233);
      $display("%x", Y234);
      $display("%x", Y235);
      $display("%x", Y236);
      $display("%x", Y237);
      $display("%x", Y238);
      $display("%x", Y239);
      $display("%x", Y240);
      $display("%x", Y241);
      $display("%x", Y242);
      $display("%x", Y243);
      $display("%x", Y244);
      $display("%x", Y245);
      $display("%x", Y246);
      $display("%x", Y247);
      $display("%x", Y248);
      $display("%x", Y249);
      $display("%x", Y250);
      $display("%x", Y251);
      $display("%x", Y252);
      $display("%x", Y253);
      $display("%x", Y254);
      $display("%x", Y255);
      $display("%x", Y256);
      $display("%x", Y257);
      $display("%x", Y258);
      $display("%x", Y259);
      $display("%x", Y260);
      $display("%x", Y261);
      $display("%x", Y262);
      $display("%x", Y263);
      $display("%x", Y264);
      $display("%x", Y265);
      $display("%x", Y266);
      $display("%x", Y267);
      $display("%x", Y268);
      $display("%x", Y269);
      $display("%x", Y270);
      $display("%x", Y271);
      $display("%x", Y272);
      $display("%x", Y273);
      $display("%x", Y274);
      $display("%x", Y275);
      $display("%x", Y276);
      $display("%x", Y277);
      $display("%x", Y278);
      $display("%x", Y279);
      $display("%x", Y280);
      $display("%x", Y281);
      $display("%x", Y282);
      $display("%x", Y283);
      $display("%x", Y284);
      $display("%x", Y285);
      $display("%x", Y286);
      $display("%x", Y287);
      $display("%x", Y288);
      $display("%x", Y289);
      $display("%x", Y290);
      $display("%x", Y291);
      $display("%x", Y292);
      $display("%x", Y293);
      $display("%x", Y294);
      $display("%x", Y295);
      $display("%x", Y296);
      $display("%x", Y297);
      $display("%x", Y298);
      $display("%x", Y299);
      $display("%x", Y300);
      $display("%x", Y301);
      $display("%x", Y302);
      $display("%x", Y303);
      $display("%x", Y304);
      $display("%x", Y305);
      $display("%x", Y306);
      $display("%x", Y307);
      $display("%x", Y308);
      $display("%x", Y309);
      $display("%x", Y310);
      $display("%x", Y311);
      $display("%x", Y312);
      $display("%x", Y313);
      $display("%x", Y314);
      $display("%x", Y315);
      $display("%x", Y316);
      $display("%x", Y317);
      $display("%x", Y318);
      $display("%x", Y319);
      $display("%x", Y320);
      $display("%x", Y321);
      $display("%x", Y322);
      $display("%x", Y323);
      $display("%x", Y324);
      $display("%x", Y325);
      $display("%x", Y326);
      $display("%x", Y327);
      $display("%x", Y328);
      $display("%x", Y329);
      $display("%x", Y330);
      $display("%x", Y331);
      $display("%x", Y332);
      $display("%x", Y333);
      $display("%x", Y334);
      $display("%x", Y335);
      $display("%x", Y336);
      $display("%x", Y337);
      $display("%x", Y338);
      $display("%x", Y339);
      $display("%x", Y340);
      $display("%x", Y341);
      $display("%x", Y342);
      $display("%x", Y343);
      $display("%x", Y344);
      $display("%x", Y345);
      $display("%x", Y346);
      $display("%x", Y347);
      $display("%x", Y348);
      $display("%x", Y349);
      $display("%x", Y350);
      $display("%x", Y351);
      $display("%x", Y352);
      $display("%x", Y353);
      $display("%x", Y354);
      $display("%x", Y355);
      $display("%x", Y356);
      $display("%x", Y357);
      $display("%x", Y358);
      $display("%x", Y359);
      $display("%x", Y360);
      $display("%x", Y361);
      $display("%x", Y362);
      $display("%x", Y363);
      $display("%x", Y364);
      $display("%x", Y365);
      $display("%x", Y366);
      $display("%x", Y367);
      $display("%x", Y368);
      $display("%x", Y369);
      $display("%x", Y370);
      $display("%x", Y371);
      $display("%x", Y372);
      $display("%x", Y373);
      $display("%x", Y374);
      $display("%x", Y375);
      $display("%x", Y376);
      $display("%x", Y377);
      $display("%x", Y378);
      $display("%x", Y379);
      $display("%x", Y380);
      $display("%x", Y381);
      $display("%x", Y382);
      $display("%x", Y383);
      $display("%x", Y384);
      $display("%x", Y385);
      $display("%x", Y386);
      $display("%x", Y387);
      $display("%x", Y388);
      $display("%x", Y389);
      $display("%x", Y390);
      $display("%x", Y391);
      $display("%x", Y392);
      $display("%x", Y393);
      $display("%x", Y394);
      $display("%x", Y395);
      $display("%x", Y396);
      $display("%x", Y397);
      $display("%x", Y398);
      $display("%x", Y399);
      $display("%x", Y400);
      $display("%x", Y401);
      $display("%x", Y402);
      $display("%x", Y403);
      $display("%x", Y404);
      $display("%x", Y405);
      $display("%x", Y406);
      $display("%x", Y407);
      $display("%x", Y408);
      $display("%x", Y409);
      $display("%x", Y410);
      $display("%x", Y411);
      $display("%x", Y412);
      $display("%x", Y413);
      $display("%x", Y414);
      $display("%x", Y415);
      $display("%x", Y416);
      $display("%x", Y417);
      $display("%x", Y418);
      $display("%x", Y419);
      $display("%x", Y420);
      $display("%x", Y421);
      $display("%x", Y422);
      $display("%x", Y423);
      $display("%x", Y424);
      $display("%x", Y425);
      $display("%x", Y426);
      $display("%x", Y427);
      $display("%x", Y428);
      $display("%x", Y429);
      $display("%x", Y430);
      $display("%x", Y431);
      $display("%x", Y432);
      $display("%x", Y433);
      $display("%x", Y434);
      $display("%x", Y435);
      $display("%x", Y436);
      $display("%x", Y437);
      $display("%x", Y438);
      $display("%x", Y439);
      $display("%x", Y440);
      $display("%x", Y441);
      $display("%x", Y442);
      $display("%x", Y443);
      $display("%x", Y444);
      $display("%x", Y445);
      $display("%x", Y446);
      $display("%x", Y447);
      $display("%x", Y448);
      $display("%x", Y449);
      $display("%x", Y450);
      $display("%x", Y451);
      $display("%x", Y452);
      $display("%x", Y453);
      $display("%x", Y454);
      $display("%x", Y455);
      $display("%x", Y456);
      $display("%x", Y457);
      $display("%x", Y458);
      $display("%x", Y459);
      $display("%x", Y460);
      $display("%x", Y461);
      $display("%x", Y462);
      $display("%x", Y463);
      $display("%x", Y464);
      $display("%x", Y465);
      $display("%x", Y466);
      $display("%x", Y467);
      $display("%x", Y468);
      $display("%x", Y469);
      $display("%x", Y470);
      $display("%x", Y471);
      $display("%x", Y472);
      $display("%x", Y473);
      $display("%x", Y474);
      $display("%x", Y475);
      $display("%x", Y476);
      $display("%x", Y477);
      $display("%x", Y478);
      $display("%x", Y479);
      $display("%x", Y480);
      $display("%x", Y481);
      $display("%x", Y482);
      $display("%x", Y483);
      $display("%x", Y484);
      $display("%x", Y485);
      $display("%x", Y486);
      $display("%x", Y487);
      $display("%x", Y488);
      $display("%x", Y489);
      $display("%x", Y490);
      $display("%x", Y491);
      $display("%x", Y492);
      $display("%x", Y493);
      $display("%x", Y494);
      $display("%x", Y495);
      $display("%x", Y496);
      $display("%x", Y497);
      $display("%x", Y498);
      $display("%x", Y499);
      $display("%x", Y500);
      $display("%x", Y501);
      $display("%x", Y502);
      $display("%x", Y503);
      $display("%x", Y504);
      $display("%x", Y505);
      $display("%x", Y506);
      $display("%x", Y507);
      $display("%x", Y508);
      $display("%x", Y509);
      $display("%x", Y510);
      $display("%x", Y511);
      $display("%x", Y512);
      $display("%x", Y513);
      $display("%x", Y514);
      $display("%x", Y515);
      $display("%x", Y516);
      $display("%x", Y517);
      $display("%x", Y518);
      $display("%x", Y519);
      $display("%x", Y520);
      $display("%x", Y521);
      $display("%x", Y522);
      $display("%x", Y523);
      $display("%x", Y524);
      $display("%x", Y525);
      $display("%x", Y526);
      $display("%x", Y527);
      $display("%x", Y528);
      $display("%x", Y529);
      $display("%x", Y530);
      $display("%x", Y531);
      $display("%x", Y532);
      $display("%x", Y533);
      $display("%x", Y534);
      $display("%x", Y535);
      $display("%x", Y536);
      $display("%x", Y537);
      $display("%x", Y538);
      $display("%x", Y539);
      $display("%x", Y540);
      $display("%x", Y541);
      $display("%x", Y542);
      $display("%x", Y543);
      $display("%x", Y544);
      $display("%x", Y545);
      $display("%x", Y546);
      $display("%x", Y547);
      $display("%x", Y548);
      $display("%x", Y549);
      $display("%x", Y550);
      $display("%x", Y551);
      $display("%x", Y552);
      $display("%x", Y553);
      $display("%x", Y554);
      $display("%x", Y555);
      $display("%x", Y556);
      $display("%x", Y557);
      $display("%x", Y558);
      $display("%x", Y559);
      $display("%x", Y560);
      $display("%x", Y561);
      $display("%x", Y562);
      $display("%x", Y563);
      $display("%x", Y564);
      $display("%x", Y565);
      $display("%x", Y566);
      $display("%x", Y567);
      $display("%x", Y568);
      $display("%x", Y569);
      $display("%x", Y570);
      $display("%x", Y571);
      $display("%x", Y572);
      $display("%x", Y573);
      $display("%x", Y574);
      $display("%x", Y575);
      $display("%x", Y576);
      $display("%x", Y577);
      $display("%x", Y578);
      $display("%x", Y579);
      $display("%x", Y580);
      $display("%x", Y581);
      $display("%x", Y582);
      $display("%x", Y583);
      $display("%x", Y584);
      $display("%x", Y585);
      $display("%x", Y586);
      $display("%x", Y587);
      $display("%x", Y588);
      $display("%x", Y589);
      $display("%x", Y590);
      $display("%x", Y591);
      $display("%x", Y592);
      $display("%x", Y593);
      $display("%x", Y594);
      $display("%x", Y595);
      $display("%x", Y596);
      $display("%x", Y597);
      $display("%x", Y598);
      $display("%x", Y599);
      $display("%x", Y600);
      $display("%x", Y601);
      $display("%x", Y602);
      $display("%x", Y603);
      $display("%x", Y604);
      $display("%x", Y605);
      $display("%x", Y606);
      $display("%x", Y607);
      $display("%x", Y608);
      $display("%x", Y609);
      $display("%x", Y610);
      $display("%x", Y611);
      $display("%x", Y612);
      $display("%x", Y613);
      $display("%x", Y614);
      $display("%x", Y615);
      $display("%x", Y616);
      $display("%x", Y617);
      $display("%x", Y618);
      $display("%x", Y619);
      $display("%x", Y620);
      $display("%x", Y621);
      $display("%x", Y622);
      $display("%x", Y623);
      $display("%x", Y624);
      $display("%x", Y625);
      $display("%x", Y626);
      $display("%x", Y627);
      $display("%x", Y628);
      $display("%x", Y629);
      $display("%x", Y630);
      $display("%x", Y631);
      $display("%x", Y632);
      $display("%x", Y633);
      $display("%x", Y634);
      $display("%x", Y635);
      $display("%x", Y636);
      $display("%x", Y637);
      $display("%x", Y638);
      $display("%x", Y639);
      $display("%x", Y640);
      $display("%x", Y641);
      $display("%x", Y642);
      $display("%x", Y643);
      $display("%x", Y644);
      $display("%x", Y645);
      $display("%x", Y646);
      $display("%x", Y647);
      $display("%x", Y648);
      $display("%x", Y649);
      $display("%x", Y650);
      $display("%x", Y651);
      $display("%x", Y652);
      $display("%x", Y653);
      $display("%x", Y654);
      $display("%x", Y655);
      $display("%x", Y656);
      $display("%x", Y657);
      $display("%x", Y658);
      $display("%x", Y659);
      $display("%x", Y660);
      $display("%x", Y661);
      $display("%x", Y662);
      $display("%x", Y663);
      $display("%x", Y664);
      $display("%x", Y665);
      $display("%x", Y666);
      $display("%x", Y667);
      $display("%x", Y668);
      $display("%x", Y669);
      $display("%x", Y670);
      $display("%x", Y671);
      $display("%x", Y672);
      $display("%x", Y673);
      $display("%x", Y674);
      $display("%x", Y675);
      $display("%x", Y676);
      $display("%x", Y677);
      $display("%x", Y678);
      $display("%x", Y679);
      $display("%x", Y680);
      $display("%x", Y681);
      $display("%x", Y682);
      $display("%x", Y683);
      $display("%x", Y684);
      $display("%x", Y685);
      $display("%x", Y686);
      $display("%x", Y687);
      $display("%x", Y688);
      $display("%x", Y689);
      $display("%x", Y690);
      $display("%x", Y691);
      $display("%x", Y692);
      $display("%x", Y693);
      $display("%x", Y694);
      $display("%x", Y695);
      $display("%x", Y696);
      $display("%x", Y697);
      $display("%x", Y698);
      $display("%x", Y699);
      $display("%x", Y700);
      $display("%x", Y701);
      $display("%x", Y702);
      $display("%x", Y703);
      $display("%x", Y704);
      $display("%x", Y705);
      $display("%x", Y706);
      $display("%x", Y707);
      $display("%x", Y708);
      $display("%x", Y709);
      $display("%x", Y710);
      $display("%x", Y711);
      $display("%x", Y712);
      $display("%x", Y713);
      $display("%x", Y714);
      $display("%x", Y715);
      $display("%x", Y716);
      $display("%x", Y717);
      $display("%x", Y718);
      $display("%x", Y719);
      $display("%x", Y720);
      $display("%x", Y721);
      $display("%x", Y722);
      $display("%x", Y723);
      $display("%x", Y724);
      $display("%x", Y725);
      $display("%x", Y726);
      $display("%x", Y727);
      $display("%x", Y728);
      $display("%x", Y729);
      $display("%x", Y730);
      $display("%x", Y731);
      $display("%x", Y732);
      $display("%x", Y733);
      $display("%x", Y734);
      $display("%x", Y735);
      $display("%x", Y736);
      $display("%x", Y737);
      $display("%x", Y738);
      $display("%x", Y739);
      $display("%x", Y740);
      $display("%x", Y741);
      $display("%x", Y742);
      $display("%x", Y743);
      $display("%x", Y744);
      $display("%x", Y745);
      $display("%x", Y746);
      $display("%x", Y747);
      $display("%x", Y748);
      $display("%x", Y749);
      $display("%x", Y750);
      $display("%x", Y751);
      $display("%x", Y752);
      $display("%x", Y753);
      $display("%x", Y754);
      $display("%x", Y755);
      $display("%x", Y756);
      $display("%x", Y757);
      $display("%x", Y758);
      $display("%x", Y759);
      $display("%x", Y760);
      $display("%x", Y761);
      $display("%x", Y762);
      $display("%x", Y763);
      $display("%x", Y764);
      $display("%x", Y765);
      $display("%x", Y766);
      $display("%x", Y767);
      $display("%x", Y768);
      $display("%x", Y769);
      $display("%x", Y770);
      $display("%x", Y771);
      $display("%x", Y772);
      $display("%x", Y773);
      $display("%x", Y774);
      $display("%x", Y775);
      $display("%x", Y776);
      $display("%x", Y777);
      $display("%x", Y778);
      $display("%x", Y779);
      $display("%x", Y780);
      $display("%x", Y781);
      $display("%x", Y782);
      $display("%x", Y783);
      $display("%x", Y784);
      $display("%x", Y785);
      $display("%x", Y786);
      $display("%x", Y787);
      $display("%x", Y788);
      $display("%x", Y789);
      $display("%x", Y790);
      $display("%x", Y791);
      $display("%x", Y792);
      $display("%x", Y793);
      $display("%x", Y794);
      $display("%x", Y795);
      $display("%x", Y796);
      $display("%x", Y797);
      $display("%x", Y798);
      $display("%x", Y799);
      $display("%x", Y800);
      $display("%x", Y801);
      $display("%x", Y802);
      $display("%x", Y803);
      $display("%x", Y804);
      $display("%x", Y805);
      $display("%x", Y806);
      $display("%x", Y807);
      $display("%x", Y808);
      $display("%x", Y809);
      $display("%x", Y810);
      $display("%x", Y811);
      $display("%x", Y812);
      $display("%x", Y813);
      $display("%x", Y814);
      $display("%x", Y815);
      $display("%x", Y816);
      $display("%x", Y817);
      $display("%x", Y818);
      $display("%x", Y819);
      $display("%x", Y820);
      $display("%x", Y821);
      $display("%x", Y822);
      $display("%x", Y823);
      $display("%x", Y824);
      $display("%x", Y825);
      $display("%x", Y826);
      $display("%x", Y827);
      $display("%x", Y828);
      $display("%x", Y829);
      $display("%x", Y830);
      $display("%x", Y831);
      $display("%x", Y832);
      $display("%x", Y833);
      $display("%x", Y834);
      $display("%x", Y835);
      $display("%x", Y836);
      $display("%x", Y837);
      $display("%x", Y838);
      $display("%x", Y839);
      $display("%x", Y840);
      $display("%x", Y841);
      $display("%x", Y842);
      $display("%x", Y843);
      $display("%x", Y844);
      $display("%x", Y845);
      $display("%x", Y846);
      $display("%x", Y847);
      $display("%x", Y848);
      $display("%x", Y849);
      $display("%x", Y850);
      $display("%x", Y851);
      $display("%x", Y852);
      $display("%x", Y853);
      $display("%x", Y854);
      $display("%x", Y855);
      $display("%x", Y856);
      $display("%x", Y857);
      $display("%x", Y858);
      $display("%x", Y859);
      $display("%x", Y860);
      $display("%x", Y861);
      $display("%x", Y862);
      $display("%x", Y863);
      $display("%x", Y864);
      $display("%x", Y865);
      $display("%x", Y866);
      $display("%x", Y867);
      $display("%x", Y868);
      $display("%x", Y869);
      $display("%x", Y870);
      $display("%x", Y871);
      $display("%x", Y872);
      $display("%x", Y873);
      $display("%x", Y874);
      $display("%x", Y875);
      $display("%x", Y876);
      $display("%x", Y877);
      $display("%x", Y878);
      $display("%x", Y879);
      $display("%x", Y880);
      $display("%x", Y881);
      $display("%x", Y882);
      $display("%x", Y883);
      $display("%x", Y884);
      $display("%x", Y885);
      $display("%x", Y886);
      $display("%x", Y887);
      $display("%x", Y888);
      $display("%x", Y889);
      $display("%x", Y890);
      $display("%x", Y891);
      $display("%x", Y892);
      $display("%x", Y893);
      $display("%x", Y894);
      $display("%x", Y895);
      $display("%x", Y896);
      $display("%x", Y897);
      $display("%x", Y898);
      $display("%x", Y899);
      $display("%x", Y900);
      $display("%x", Y901);
      $display("%x", Y902);
      $display("%x", Y903);
      $display("%x", Y904);
      $display("%x", Y905);
      $display("%x", Y906);
      $display("%x", Y907);
      $display("%x", Y908);
      $display("%x", Y909);
      $display("%x", Y910);
      $display("%x", Y911);
      $display("%x", Y912);
      $display("%x", Y913);
      $display("%x", Y914);
      $display("%x", Y915);
      $display("%x", Y916);
      $display("%x", Y917);
      $display("%x", Y918);
      $display("%x", Y919);
      $display("%x", Y920);
      $display("%x", Y921);
      $display("%x", Y922);
      $display("%x", Y923);
      $display("%x", Y924);
      $display("%x", Y925);
      $display("%x", Y926);
      $display("%x", Y927);
      $display("%x", Y928);
      $display("%x", Y929);
      $display("%x", Y930);
      $display("%x", Y931);
      $display("%x", Y932);
      $display("%x", Y933);
      $display("%x", Y934);
      $display("%x", Y935);
      $display("%x", Y936);
      $display("%x", Y937);
      $display("%x", Y938);
      $display("%x", Y939);
      $display("%x", Y940);
      $display("%x", Y941);
      $display("%x", Y942);
      $display("%x", Y943);
      $display("%x", Y944);
      $display("%x", Y945);
      $display("%x", Y946);
      $display("%x", Y947);
      $display("%x", Y948);
      $display("%x", Y949);
      $display("%x", Y950);
      $display("%x", Y951);
      $display("%x", Y952);
      $display("%x", Y953);
      $display("%x", Y954);
      $display("%x", Y955);
      $display("%x", Y956);
      $display("%x", Y957);
      $display("%x", Y958);
      $display("%x", Y959);
      $display("%x", Y960);
      $display("%x", Y961);
      $display("%x", Y962);
      $display("%x", Y963);
      $display("%x", Y964);
      $display("%x", Y965);
      $display("%x", Y966);
      $display("%x", Y967);
      $display("%x", Y968);
      $display("%x", Y969);
      $display("%x", Y970);
      $display("%x", Y971);
      $display("%x", Y972);
      $display("%x", Y973);
      $display("%x", Y974);
      $display("%x", Y975);
      $display("%x", Y976);
      $display("%x", Y977);
      $display("%x", Y978);
      $display("%x", Y979);
      $display("%x", Y980);
      $display("%x", Y981);
      $display("%x", Y982);
      $display("%x", Y983);
      $display("%x", Y984);
      $display("%x", Y985);
      $display("%x", Y986);
      $display("%x", Y987);
      $display("%x", Y988);
      $display("%x", Y989);
      $display("%x", Y990);
      $display("%x", Y991);
      $display("%x", Y992);
      $display("%x", Y993);
      $display("%x", Y994);
      $display("%x", Y995);
      $display("%x", Y996);
      $display("%x", Y997);
      $display("%x", Y998);
      $display("%x", Y999);
      $display("%x", Y1000);
      $display("%x", Y1001);
      $display("%x", Y1002);
      $display("%x", Y1003);
      $display("%x", Y1004);
      $display("%x", Y1005);
      $display("%x", Y1006);
      $display("%x", Y1007);
      $display("%x", Y1008);
      $display("%x", Y1009);
      $display("%x", Y1010);
      $display("%x", Y1011);
      $display("%x", Y1012);
      $display("%x", Y1013);
      $display("%x", Y1014);
      $display("%x", Y1015);
      $display("%x", Y1016);
      $display("%x", Y1017);
      $display("%x", Y1018);
      $display("%x", Y1019);
      $display("%x", Y1020);
      $display("%x", Y1021);
      $display("%x", Y1022);
      $display("%x", Y1023);
      $finish;
   end
endmodule
